`default_nettype none

(* blackbox *)
module fa16b_rev (
    inout  wire vss,
    inout  wire vdd,
    inout wire c15,
    inout wire c15_not,
    inout  wire c0_f_not,
    inout  wire a0_f,
    inout  wire c0_f,
    inout  wire b0,
    inout  wire a0_f_not,
    inout  wire b1_not,
    inout  wire b0_not,
    inout  wire b1,
    inout  wire a1_not,
    inout  wire b2_not,
    inout  wire a1,
    inout  wire b2,
    inout  wire a2_not,
    inout  wire b3_not,
    inout  wire a2,
    inout  wire b3,
    inout  wire a3_not,
    inout  wire b4_not,
    inout  wire a3,
    inout  wire b4,
    inout  wire a4_not,
    inout  wire b5_not,
    inout  wire a4,
    inout  wire b5,
    inout  wire a5_not,
    inout  wire b6_not,
    inout  wire a5,
    inout  wire b6,
    inout  wire a6_not,
    inout  wire b7_not,
    inout  wire a6,
    inout  wire b7,
    inout  wire a7_not,
    inout  wire a7,
    inout  wire a7_b,
    inout wire s7,
    inout  wire a7_not_b,
    inout wire s7_not,
    inout  wire a6_b,
    inout wire s6,
    inout  wire a6_not_b,
    inout wire s6_not,
    inout  wire a5_b,
    inout wire s5,
    inout  wire a5_not_b,
    inout wire s5_not,
    inout  wire a4_b,
    inout wire s4,
    inout  wire a4_not_b,
    inout wire s4_not,
    inout  wire a3_b,
    inout wire s3,
    inout  wire a3_not_b,
    inout wire s3_not,
    inout  wire a2_b,
    inout wire s2,
    inout  wire a2_not_b,
    inout wire s2_not,
    inout  wire a1_b,
    inout wire s1,
    inout  wire a1_not_b,
    inout wire s1_not,
    inout  wire a0_b,
    inout wire s0,
    inout  wire a0_not_b,
    inout wire s0_not,
    inout  wire c0_b,
    inout  wire c0_not_b,
    inout  wire b8_not,
    inout  wire a8_not,
    inout  wire b8,
    inout  wire a8,
    inout  wire b9_not,
    inout  wire a9_not,
    inout  wire b9,
    inout  wire a9,
    inout  wire b10_not,
    inout  wire a10_not,
    inout  wire b10,
    inout  wire a10,
    inout  wire b11_not,
    inout  wire a11_not,
    inout  wire b11,
    inout  wire a11,
    inout  wire b12_not,
    inout  wire a12_not,
    inout  wire b12,
    inout  wire a12,
    inout  wire b13_not,
    inout  wire a13_not,
    inout  wire b13,
    inout  wire a13,
    inout  wire b14_not,
    inout  wire a14_not,
    inout  wire b14,
    inout  wire a14,
    inout  wire b15_not,
    inout  wire a15_not,
    inout  wire b15,
    inout  wire a15,
    inout  wire a15_b,
    inout wire s15,
    inout wire s15_not,
    inout  wire a14_b,
    inout wire s14,
    inout  wire a14_not_b,
    inout wire s14_not,
    inout  wire a13_b,
    inout wire s13,
    inout  wire a13_not_b,
    inout wire s13_not,
    inout  wire a12_b,
    inout wire s12,
    inout  wire a12_not_b,
    inout wire s12_not,
    inout  wire a11_b,
    inout wire s11,
    inout  wire a11_not_b,
    inout wire s11_not,
    inout  wire a10_b,
    inout wire s10,
    inout  wire a10_not_b,
    inout wire s10_not,
    inout  wire a9_b,
    inout wire s9,
    inout  wire a9_not_b,
    inout wire s9_not,
    inout  wire a8_b,
    inout wire s8,
    inout  wire a8_not_b,
    inout wire s8_not,
    inout  wire a15_not_b,
    inout wire z_not,
    inout wire z
);

endmodule
