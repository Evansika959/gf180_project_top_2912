`default_nettype none

module fa16_rev_wrapped (
    `ifdef USE_POWER_PINS
    inout  wire vdd,
    inout  wire vss,
    `endif

    // Input ports
    input  wire [15:0] a,
    input  wire [15:0] a_not,
    input  wire [15:0] b,
    input  wire [15:0] b_not,
    input  wire        c0_f,
    input  wire        c0_f_not,
    
    
    // Output ports
    output wire [15:0] s,
    output wire [15:0] s_not,
    output wire [15:0] a_b,
    output wire [15:0] a_not_b,
    output wire        c15,
    output wire        c15_not,
    output wire        c0_b,
    output wire        c0_not_b,
    output wire        z,
    output wire        z_not
);

    // Power handling
    `ifndef USE_POWER_PINS
    wire vdd = 1'b1;
    wire vss = 1'b0;
    `endif

    

    wire a0_f;
    wire a0_f_not;

    assign a0_f     = 1'b0;
    assign a0_f_not = 1'b1;

    (* keep *)
    fa16b_rev u_fa16b_rev (
        .vss         (vss),
        .vdd         (vdd),
        .c15         (c15),
        .c15_not     (c15_not),
        .c0_f_not    (c0_f_not),
        .a0_f        (a0_f),
        .c0_f        (c0_f),
        .b0          (b[0]),
        .a0_f_not    (a0_f_not),
        .b1_not      (b_not[1]),
        .b0_not      (b_not[0]),
        .b1          (b[1]),
        .a1_not      (a_not[1]),
        .b2_not      (b_not[2]),
        .a1          (a[1]),
        .b2          (b[2]),
        .a2_not      (a_not[2]),
        .b3_not      (b_not[3]),
        .a2          (a[2]),
        .b3          (b[3]),
        .a3_not      (a_not[3]),
        .b4_not      (b_not[4]),
        .a3          (a[3]),
        .b4          (b[4]),
        .a4_not      (a_not[4]),
        .b5_not      (b_not[5]),
        .a4          (a[4]),
        .b5          (b[5]),
        .a5_not      (a_not[5]),
        .b6_not      (b_not[6]),
        .a5          (a[5]),
        .b6          (b[6]),
        .a6_not      (a_not[6]),
        .b7_not      (b_not[7]),
        .a6          (a[6]),
        .b7          (b[7]),
        .a7_not      (a_not[7]),
        .a7          (a[7]),
    .a7_b        (a_b[7]),
    .s7          (s[7]),
    .a7_not_b    (a_not_b[7]),
    .s7_not      (s_not[7]),
    .a6_b        (a_b[6]),
    .s6          (s[6]),
    .a6_not_b    (a_not_b[6]),
    .s6_not      (s_not[6]),
    .a5_b        (a_b[5]),
    .s5          (s[5]),
    .a5_not_b    (a_not_b[5]),
    .s5_not      (s_not[5]),
    .a4_b        (a_b[4]),
    .s4          (s[4]),
    .a4_not_b    (a_not_b[4]),
    .s4_not      (s_not[4]),
    .a3_b        (a_b[3]),
    .s3          (s[3]),
    .a3_not_b    (a_not_b[3]),
    .s3_not      (s_not[3]),
    .a2_b        (a_b[2]),
    .s2          (s[2]),
    .a2_not_b    (a_not_b[2]),
    .s2_not      (s_not[2]),
    .a1_b        (a_b[1]),
    .s1          (s[1]),
    .a1_not_b    (a_not_b[1]),
    .s1_not      (s_not[1]),
    .a0_b        (a_b[0]),
    .s0          (s[0]),
    .a0_not_b    (a_not_b[0]),
    .s0_not      (s_not[0]),
        .c0_b        (c0_b),
        .c0_not_b    (c0_not_b),
        .b8_not      (b_not[8]),
        .a8_not      (a_not[8]),
        .b8          (b[8]),
        .a8          (a[8]),
        .b9_not      (b_not[9]),
        .a9_not      (a_not[9]),
        .b9          (b[9]),
        .a9          (a[9]),
        .b10_not     (b_not[10]),
        .a10_not     (a_not[10]),
        .b10         (b[10]),
        .a10         (a[10]),
        .b11_not     (b_not[11]),
        .a11_not     (a_not[11]),
        .b11         (b[11]),
        .a11         (a[11]),
        .b12_not     (b_not[12]),
        .a12_not     (a_not[12]),
        .b12         (b[12]),
        .a12         (a[12]),
        .b13_not     (b_not[13]),
        .a13_not     (a_not[13]),
        .b13         (b[13]),
        .a13         (a[13]),
        .b14_not     (b_not[14]),
        .a14_not     (a_not[14]),
        .b14         (b[14]),
        .a14         (a[14]),
        .b15_not     (b_not[15]),
        .a15_not     (a_not[15]),
        .b15         (b[15]),
        .a15         (a[15]),
    .a15_b       (a_b[15]),
    .s15         (s[15]),
    .s15_not     (s_not[15]),
    .a14_b       (a_b[14]),
    .s14         (s[14]),
    .a14_not_b   (a_not_b[14]),
    .s14_not     (s_not[14]),
    .a13_b       (a_b[13]),
    .s13         (s[13]),
    .a13_not_b   (a_not_b[13]),
    .s13_not     (s_not[13]),
    .a12_b       (a_b[12]),
    .s12         (s[12]),
    .a12_not_b   (a_not_b[12]),
    .s12_not     (s_not[12]),
    .a11_b       (a_b[11]),
    .s11         (s[11]),
    .a11_not_b   (a_not_b[11]),
    .s11_not     (s_not[11]),
    .a10_b       (a_b[10]),
    .s10         (s[10]),
    .a10_not_b   (a_not_b[10]),
    .s10_not     (s_not[10]),
    .a9_b        (a_b[9]),
    .s9          (s[9]),
    .a9_not_b    (a_not_b[9]),
    .s9_not      (s_not[9]),
    .a8_b        (a_b[8]),
    .s8          (s[8]),
    .a8_not_b    (a_not_b[8]),
    .s8_not      (s_not[8]),
        .a15_not_b   (a_not_b[15]),
        .z_not       (z_not),
        .z           (z)
    );

endmodule