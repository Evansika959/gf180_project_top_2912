VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO 8b_mult
  CLASS BLOCK ;
  FOREIGN 8b_mult ;
  ORIGIN 106.705 -0.235 ;
  SIZE 1422.930 BY 204.320 ;
  PIN b6_q0
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT 927.535 204.205 929.155 204.530 ;
        RECT 952.410 168.220 952.790 168.600 ;
        RECT 973.910 168.220 974.290 168.600 ;
        RECT 949.265 165.875 967.935 165.885 ;
        RECT 928.350 165.565 975.920 165.875 ;
        RECT 928.350 165.550 949.560 165.565 ;
        RECT 960.410 163.105 960.790 163.110 ;
        RECT 957.930 162.740 960.795 163.105 ;
        RECT 965.910 163.085 966.290 163.110 ;
        RECT 965.895 162.765 968.040 163.085 ;
        RECT 960.410 162.730 960.790 162.740 ;
        RECT 965.910 162.730 966.290 162.765 ;
        RECT 952.325 148.505 952.705 148.885 ;
        RECT 973.825 148.505 974.205 148.885 ;
        RECT 928.370 146.170 949.390 146.180 ;
        RECT 928.370 146.160 967.850 146.170 ;
        RECT 928.370 145.855 975.835 146.160 ;
        RECT 949.180 145.850 975.835 145.855 ;
        RECT 960.325 143.390 960.705 143.395 ;
        RECT 957.845 143.025 960.710 143.390 ;
        RECT 965.825 143.370 966.205 143.395 ;
        RECT 965.810 143.050 967.955 143.370 ;
        RECT 960.325 143.015 960.705 143.025 ;
        RECT 965.825 143.015 966.205 143.050 ;
        RECT 952.385 128.700 952.765 129.080 ;
        RECT 973.885 128.700 974.265 129.080 ;
        RECT 928.320 126.365 949.600 126.370 ;
        RECT 928.320 126.355 967.910 126.365 ;
        RECT 928.320 126.045 975.895 126.355 ;
        RECT 960.385 123.585 960.765 123.590 ;
        RECT 957.905 123.220 960.770 123.585 ;
        RECT 965.885 123.565 966.265 123.590 ;
        RECT 965.870 123.245 968.015 123.565 ;
        RECT 960.385 123.210 960.765 123.220 ;
        RECT 965.885 123.210 966.265 123.245 ;
        RECT 952.315 108.930 952.695 109.310 ;
        RECT 973.815 108.930 974.195 109.310 ;
        RECT 928.325 106.595 949.370 106.610 ;
        RECT 928.325 106.585 967.840 106.595 ;
        RECT 928.325 106.285 975.825 106.585 ;
        RECT 949.170 106.275 975.825 106.285 ;
        RECT 960.315 103.815 960.695 103.820 ;
        RECT 957.835 103.450 960.700 103.815 ;
        RECT 965.815 103.795 966.195 103.820 ;
        RECT 965.800 103.475 967.945 103.795 ;
        RECT 960.315 103.440 960.695 103.450 ;
        RECT 965.815 103.440 966.195 103.475 ;
        RECT 952.345 89.205 952.725 89.585 ;
        RECT 973.845 89.205 974.225 89.585 ;
        RECT 928.310 86.870 949.390 86.875 ;
        RECT 928.310 86.860 967.870 86.870 ;
        RECT 928.310 86.550 975.855 86.860 ;
        RECT 960.345 84.090 960.725 84.095 ;
        RECT 957.865 83.725 960.730 84.090 ;
        RECT 965.845 84.070 966.225 84.095 ;
        RECT 965.830 83.750 967.975 84.070 ;
        RECT 960.345 83.715 960.725 83.725 ;
        RECT 965.845 83.715 966.225 83.750 ;
        RECT 952.275 69.375 952.655 69.755 ;
        RECT 973.775 69.375 974.155 69.755 ;
        RECT 928.295 67.030 967.800 67.040 ;
        RECT 928.295 66.720 975.785 67.030 ;
        RECT 928.295 66.715 949.315 66.720 ;
        RECT 960.275 64.260 960.655 64.265 ;
        RECT 957.795 63.895 960.660 64.260 ;
        RECT 965.775 64.240 966.155 64.265 ;
        RECT 965.760 63.920 967.905 64.240 ;
        RECT 960.275 63.885 960.655 63.895 ;
        RECT 965.775 63.885 966.155 63.920 ;
        RECT 952.345 49.655 952.725 50.035 ;
        RECT 973.845 49.655 974.225 50.035 ;
        RECT 928.405 47.320 949.455 47.330 ;
        RECT 928.405 47.310 967.870 47.320 ;
        RECT 928.405 47.005 975.855 47.310 ;
        RECT 949.200 47.000 975.855 47.005 ;
        RECT 960.345 44.540 960.725 44.545 ;
        RECT 957.865 44.175 960.730 44.540 ;
        RECT 965.845 44.520 966.225 44.545 ;
        RECT 965.830 44.200 967.975 44.520 ;
        RECT 960.345 44.165 960.725 44.175 ;
        RECT 965.845 44.165 966.225 44.200 ;
        RECT 952.320 29.925 952.700 30.305 ;
        RECT 973.820 29.925 974.200 30.305 ;
        RECT 949.175 27.585 967.845 27.590 ;
        RECT 928.340 27.580 967.845 27.585 ;
        RECT 928.340 27.270 975.830 27.580 ;
        RECT 928.340 27.260 949.320 27.270 ;
        RECT 960.320 24.810 960.700 24.815 ;
        RECT 957.840 24.445 960.705 24.810 ;
        RECT 965.820 24.790 966.200 24.815 ;
        RECT 965.805 24.470 967.950 24.790 ;
        RECT 960.320 24.435 960.700 24.445 ;
        RECT 965.820 24.435 966.200 24.470 ;
      LAYER Metal2 ;
        RECT 928.560 17.835 928.955 204.530 ;
        RECT 952.360 165.565 952.810 168.555 ;
        RECT 958.085 162.555 958.490 165.885 ;
        RECT 967.520 162.610 967.970 165.885 ;
        RECT 973.875 165.565 974.325 168.575 ;
        RECT 952.275 145.850 952.725 148.840 ;
        RECT 958.000 142.840 958.405 146.170 ;
        RECT 967.435 142.895 967.885 146.170 ;
        RECT 973.790 145.850 974.240 148.860 ;
        RECT 952.335 126.045 952.785 129.035 ;
        RECT 958.060 123.035 958.465 126.365 ;
        RECT 967.495 123.090 967.945 126.365 ;
        RECT 973.850 126.045 974.300 129.055 ;
        RECT 952.265 106.275 952.715 109.265 ;
        RECT 957.990 103.265 958.395 106.595 ;
        RECT 967.425 103.320 967.875 106.595 ;
        RECT 973.780 106.275 974.230 109.285 ;
        RECT 952.295 86.550 952.745 89.540 ;
        RECT 958.020 83.540 958.425 86.870 ;
        RECT 967.455 83.595 967.905 86.870 ;
        RECT 973.810 86.550 974.260 89.560 ;
        RECT 952.225 66.720 952.675 69.710 ;
        RECT 957.950 63.710 958.355 67.040 ;
        RECT 967.385 63.765 967.835 67.040 ;
        RECT 973.740 66.720 974.190 69.730 ;
        RECT 952.295 47.000 952.745 49.990 ;
        RECT 958.020 43.990 958.425 47.320 ;
        RECT 967.455 44.045 967.905 47.320 ;
        RECT 973.810 47.000 974.260 50.010 ;
        RECT 952.270 27.270 952.720 30.260 ;
        RECT 957.995 24.260 958.400 27.590 ;
        RECT 967.430 24.315 967.880 27.590 ;
        RECT 973.785 27.270 974.235 30.280 ;
    END
  END b6_q0
  PIN b6_q0_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT 927.520 203.630 930.080 203.935 ;
        RECT 956.410 168.220 956.790 168.600 ;
        RECT 969.910 168.220 970.290 168.600 ;
        RECT 949.265 164.885 975.920 164.895 ;
        RECT 929.510 164.625 975.920 164.885 ;
        RECT 929.510 164.615 949.505 164.625 ;
        RECT 952.410 163.075 952.790 163.110 ;
        RECT 973.910 163.090 974.290 163.110 ;
        RECT 952.145 162.765 955.155 163.075 ;
        RECT 971.445 162.770 974.355 163.090 ;
        RECT 952.410 162.730 952.790 162.765 ;
        RECT 973.910 162.730 974.290 162.770 ;
        RECT 956.325 148.505 956.705 148.885 ;
        RECT 969.825 148.505 970.205 148.885 ;
        RECT 929.530 145.180 949.335 145.190 ;
        RECT 929.530 144.920 975.835 145.180 ;
        RECT 949.180 144.910 975.835 144.920 ;
        RECT 952.325 143.360 952.705 143.395 ;
        RECT 973.825 143.375 974.205 143.395 ;
        RECT 952.060 143.050 955.070 143.360 ;
        RECT 971.360 143.055 974.270 143.375 ;
        RECT 952.325 143.015 952.705 143.050 ;
        RECT 973.825 143.015 974.205 143.055 ;
        RECT 956.385 128.700 956.765 129.080 ;
        RECT 969.885 128.700 970.265 129.080 ;
        RECT 929.480 125.375 949.565 125.380 ;
        RECT 929.480 125.110 975.895 125.375 ;
        RECT 949.240 125.105 975.895 125.110 ;
        RECT 952.385 123.555 952.765 123.590 ;
        RECT 973.885 123.570 974.265 123.590 ;
        RECT 952.120 123.245 955.130 123.555 ;
        RECT 971.420 123.250 974.330 123.570 ;
        RECT 952.385 123.210 952.765 123.245 ;
        RECT 973.885 123.210 974.265 123.250 ;
        RECT 956.315 108.930 956.695 109.310 ;
        RECT 969.815 108.930 970.195 109.310 ;
        RECT 929.485 105.605 949.390 105.620 ;
        RECT 929.485 105.350 975.825 105.605 ;
        RECT 949.170 105.335 975.825 105.350 ;
        RECT 952.315 103.785 952.695 103.820 ;
        RECT 973.815 103.800 974.195 103.820 ;
        RECT 952.050 103.475 955.060 103.785 ;
        RECT 971.350 103.480 974.260 103.800 ;
        RECT 952.315 103.440 952.695 103.475 ;
        RECT 973.815 103.440 974.195 103.480 ;
        RECT 956.345 89.205 956.725 89.585 ;
        RECT 969.845 89.205 970.225 89.585 ;
        RECT 929.470 85.880 949.445 85.885 ;
        RECT 929.470 85.615 975.855 85.880 ;
        RECT 949.200 85.610 975.855 85.615 ;
        RECT 952.345 84.060 952.725 84.095 ;
        RECT 973.845 84.075 974.225 84.095 ;
        RECT 952.080 83.750 955.090 84.060 ;
        RECT 971.380 83.755 974.290 84.075 ;
        RECT 952.345 83.715 952.725 83.750 ;
        RECT 973.845 83.715 974.225 83.755 ;
        RECT 956.275 69.375 956.655 69.755 ;
        RECT 969.775 69.375 970.155 69.755 ;
        RECT 929.450 65.780 975.785 66.050 ;
        RECT 952.275 64.230 952.655 64.265 ;
        RECT 973.775 64.245 974.155 64.265 ;
        RECT 952.010 63.920 955.020 64.230 ;
        RECT 971.310 63.925 974.220 64.245 ;
        RECT 952.275 63.885 952.655 63.920 ;
        RECT 973.775 63.885 974.155 63.925 ;
        RECT 956.345 49.655 956.725 50.035 ;
        RECT 969.845 49.655 970.225 50.035 ;
        RECT 929.565 46.330 949.455 46.340 ;
        RECT 929.565 46.070 975.855 46.330 ;
        RECT 949.200 46.060 975.855 46.070 ;
        RECT 952.345 44.510 952.725 44.545 ;
        RECT 973.845 44.525 974.225 44.545 ;
        RECT 952.080 44.200 955.090 44.510 ;
        RECT 971.380 44.205 974.290 44.525 ;
        RECT 952.345 44.165 952.725 44.200 ;
        RECT 973.845 44.165 974.225 44.205 ;
        RECT 956.320 29.925 956.700 30.305 ;
        RECT 969.820 29.925 970.200 30.305 ;
        RECT 949.175 26.595 975.830 26.600 ;
        RECT 929.500 26.330 975.830 26.595 ;
        RECT 929.500 26.325 949.400 26.330 ;
        RECT 952.320 24.780 952.700 24.815 ;
        RECT 973.820 24.795 974.200 24.815 ;
        RECT 952.055 24.470 955.065 24.780 ;
        RECT 971.355 24.475 974.265 24.795 ;
        RECT 952.320 24.435 952.700 24.470 ;
        RECT 973.820 24.435 974.200 24.475 ;
      LAYER Metal2 ;
        RECT 929.665 17.920 930.005 204.520 ;
        RECT 954.760 162.580 955.055 164.950 ;
        RECT 956.370 164.625 956.820 168.590 ;
        RECT 969.900 164.625 970.300 168.565 ;
        RECT 971.550 162.615 971.965 165.005 ;
        RECT 954.675 142.865 954.970 145.235 ;
        RECT 956.285 144.910 956.735 148.875 ;
        RECT 969.815 144.910 970.215 148.850 ;
        RECT 971.465 142.900 971.880 145.290 ;
        RECT 954.735 123.060 955.030 125.430 ;
        RECT 956.345 125.105 956.795 129.070 ;
        RECT 969.875 125.105 970.275 129.045 ;
        RECT 971.525 123.095 971.940 125.485 ;
        RECT 954.665 103.290 954.960 105.660 ;
        RECT 956.275 105.335 956.725 109.300 ;
        RECT 969.805 105.335 970.205 109.275 ;
        RECT 971.455 103.325 971.870 105.715 ;
        RECT 954.695 83.565 954.990 85.935 ;
        RECT 956.305 85.610 956.755 89.575 ;
        RECT 969.835 85.610 970.235 89.550 ;
        RECT 971.485 83.600 971.900 85.990 ;
        RECT 954.625 63.735 954.920 66.105 ;
        RECT 956.235 65.780 956.685 69.745 ;
        RECT 969.765 65.780 970.165 69.720 ;
        RECT 971.415 63.770 971.830 66.160 ;
        RECT 954.695 44.015 954.990 46.385 ;
        RECT 956.305 46.060 956.755 50.025 ;
        RECT 969.835 46.060 970.235 50.000 ;
        RECT 971.485 44.050 971.900 46.440 ;
        RECT 954.670 24.285 954.965 26.655 ;
        RECT 956.280 26.330 956.730 30.295 ;
        RECT 969.810 26.330 970.210 30.270 ;
        RECT 971.460 24.320 971.875 26.710 ;
    END
  END b6_q0_not
  PIN b6_p0_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.645 202.485 1143.735 202.815 ;
        RECT -21.310 188.205 -20.930 188.250 ;
        RECT -15.810 188.205 -15.430 188.250 ;
        RECT -21.360 187.890 -15.425 188.205 ;
        RECT -21.310 187.870 -20.930 187.890 ;
        RECT -15.810 187.870 -15.430 187.890 ;
        RECT -29.310 180.380 -28.220 180.760 ;
        RECT -7.810 180.715 -7.430 180.760 ;
        RECT -8.545 180.415 -7.235 180.715 ;
        RECT -7.810 180.380 -7.430 180.415 ;
        RECT -50.095 179.870 -32.075 179.955 ;
        RECT -50.095 179.605 -5.800 179.870 ;
        RECT -32.455 179.520 -5.800 179.605 ;
        RECT 174.950 168.560 175.330 168.605 ;
        RECT 180.450 168.560 180.830 168.605 ;
        RECT 567.660 168.565 568.040 168.610 ;
        RECT 573.160 168.565 573.540 168.610 ;
        RECT 764.025 168.570 764.405 168.615 ;
        RECT 769.525 168.570 769.905 168.615 ;
        RECT -71.545 168.470 -71.165 168.515 ;
        RECT -66.045 168.470 -65.665 168.515 ;
        RECT -71.595 168.155 -65.660 168.470 ;
        RECT 174.900 168.245 180.835 168.560 ;
        RECT 371.340 168.520 371.720 168.565 ;
        RECT 376.840 168.520 377.220 168.565 ;
        RECT 174.950 168.225 175.330 168.245 ;
        RECT 180.450 168.225 180.830 168.245 ;
        RECT 371.290 168.205 377.225 168.520 ;
        RECT 567.610 168.250 573.545 168.565 ;
        RECT 763.975 168.255 769.910 168.570 ;
        RECT 960.410 168.555 960.790 168.600 ;
        RECT 965.910 168.555 966.290 168.600 ;
        RECT 1156.735 168.560 1157.115 168.605 ;
        RECT 1162.235 168.560 1162.615 168.605 ;
        RECT 567.660 168.230 568.040 168.250 ;
        RECT 573.160 168.230 573.540 168.250 ;
        RECT 764.025 168.235 764.405 168.255 ;
        RECT 769.525 168.235 769.905 168.255 ;
        RECT 960.360 168.240 966.295 168.555 ;
        RECT 1156.685 168.245 1162.620 168.560 ;
        RECT 960.410 168.220 960.790 168.240 ;
        RECT 965.910 168.220 966.290 168.240 ;
        RECT 1156.735 168.225 1157.115 168.245 ;
        RECT 1162.235 168.225 1162.615 168.245 ;
        RECT 371.340 168.185 371.720 168.205 ;
        RECT 376.840 168.185 377.220 168.205 ;
        RECT -71.545 168.135 -71.165 168.155 ;
        RECT -66.045 168.135 -65.665 168.155 ;
        RECT -79.545 160.645 -78.455 161.025 ;
        RECT -58.045 160.980 -57.665 161.025 ;
        RECT -58.780 160.680 -57.470 160.980 ;
        RECT 166.950 160.735 168.040 161.115 ;
        RECT 188.450 161.070 188.830 161.115 ;
        RECT 187.715 160.770 189.025 161.070 ;
        RECT 188.450 160.735 188.830 160.770 ;
        RECT 363.340 160.695 364.430 161.075 ;
        RECT 384.840 161.030 385.220 161.075 ;
        RECT 384.105 160.730 385.415 161.030 ;
        RECT 559.660 160.740 560.750 161.120 ;
        RECT 581.160 161.075 581.540 161.120 ;
        RECT 580.425 160.775 581.735 161.075 ;
        RECT 581.160 160.740 581.540 160.775 ;
        RECT 756.025 160.745 757.115 161.125 ;
        RECT 777.525 161.080 777.905 161.125 ;
        RECT 776.790 160.780 778.100 161.080 ;
        RECT 777.525 160.745 777.905 160.780 ;
        RECT 952.410 160.730 953.500 161.110 ;
        RECT 973.910 161.065 974.290 161.110 ;
        RECT 973.175 160.765 974.485 161.065 ;
        RECT 973.910 160.730 974.290 160.765 ;
        RECT 1148.735 160.735 1149.825 161.115 ;
        RECT 1170.235 161.070 1170.615 161.115 ;
        RECT 1169.500 160.770 1170.810 161.070 ;
        RECT 1170.235 160.735 1170.615 160.770 ;
        RECT 384.840 160.695 385.220 160.730 ;
        RECT -58.045 160.645 -57.665 160.680 ;
        RECT 163.805 160.215 190.460 160.225 ;
        RECT 556.515 160.220 583.170 160.230 ;
        RECT 752.880 160.225 779.535 160.235 ;
        RECT -99.860 159.785 -56.035 160.135 ;
        RECT 146.080 159.875 190.460 160.215 ;
        RECT 360.195 160.175 386.850 160.185 ;
        RECT 146.080 159.865 164.100 159.875 ;
        RECT 342.470 159.835 386.850 160.175 ;
        RECT 538.790 159.880 583.170 160.220 ;
        RECT 735.155 159.885 779.535 160.225 ;
        RECT 949.265 160.210 975.920 160.220 ;
        RECT 1145.590 160.215 1172.245 160.225 ;
        RECT 538.790 159.870 556.810 159.880 ;
        RECT 735.155 159.875 753.175 159.885 ;
        RECT 931.540 159.870 975.920 160.210 ;
        RECT 1127.865 159.875 1172.245 160.215 ;
        RECT 931.540 159.860 949.560 159.870 ;
        RECT 1127.865 159.865 1145.885 159.875 ;
        RECT 342.470 159.825 360.490 159.835 ;
      LAYER Metal2 ;
        RECT -99.690 18.040 -99.405 204.535 ;
        RECT -78.930 159.785 -78.550 161.160 ;
        RECT -69.220 159.495 -68.850 168.595 ;
        RECT -58.675 159.700 -58.340 161.050 ;
        RECT -49.930 17.850 -49.645 204.500 ;
        RECT -28.695 179.520 -28.315 180.895 ;
        RECT -18.985 179.230 -18.615 188.330 ;
        RECT -8.440 179.435 -8.105 180.785 ;
        RECT 146.240 17.860 146.525 204.510 ;
        RECT 167.565 159.875 167.945 161.250 ;
        RECT 177.275 159.585 177.645 168.685 ;
        RECT 187.820 159.790 188.155 161.140 ;
        RECT 342.630 17.820 342.915 204.470 ;
        RECT 363.955 159.835 364.335 161.210 ;
        RECT 373.665 159.545 374.035 168.645 ;
        RECT 384.210 159.750 384.545 161.100 ;
        RECT 538.950 17.865 539.235 204.515 ;
        RECT 560.275 159.880 560.655 161.255 ;
        RECT 569.985 159.590 570.355 168.690 ;
        RECT 580.530 159.795 580.865 161.145 ;
        RECT 735.315 17.870 735.600 204.520 ;
        RECT 756.640 159.885 757.020 161.260 ;
        RECT 766.350 159.595 766.720 168.695 ;
        RECT 776.895 159.800 777.230 161.150 ;
        RECT 931.700 17.855 931.985 204.505 ;
        RECT 953.025 159.870 953.405 161.245 ;
        RECT 962.735 159.580 963.105 168.680 ;
        RECT 973.280 159.785 973.615 161.135 ;
        RECT 1128.025 17.860 1128.310 204.510 ;
        RECT 1149.350 159.875 1149.730 161.250 ;
        RECT 1159.060 159.585 1159.430 168.685 ;
        RECT 1169.605 159.790 1169.940 161.140 ;
    END
  END b6_p0_not
  PIN b6_p0
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.665 203.075 1143.740 203.360 ;
        RECT -51.060 192.065 -32.155 192.150 ;
        RECT -51.060 191.865 -5.800 192.065 ;
        RECT -32.455 191.780 -5.800 191.865 ;
        RECT -7.810 190.615 -7.430 190.650 ;
        RECT -29.310 190.510 -28.930 190.550 ;
        RECT -29.380 190.205 -26.545 190.510 ;
        RECT -10.565 190.305 -7.430 190.615 ;
        RECT -7.810 190.270 -7.430 190.305 ;
        RECT -29.310 190.170 -28.930 190.205 ;
        RECT -25.310 182.380 -24.220 182.760 ;
        RECT -12.765 182.380 -11.430 182.760 ;
        RECT -24.825 180.385 -11.975 180.720 ;
        RECT 163.805 172.410 190.460 172.420 ;
        RECT 556.515 172.415 583.170 172.425 ;
        RECT 752.880 172.420 779.535 172.430 ;
        RECT -100.825 172.045 -56.035 172.330 ;
        RECT 145.115 172.135 190.460 172.410 ;
        RECT 360.195 172.370 386.850 172.380 ;
        RECT 145.115 172.125 164.020 172.135 ;
        RECT 341.505 172.095 386.850 172.370 ;
        RECT 537.825 172.140 583.170 172.415 ;
        RECT 734.190 172.145 779.535 172.420 ;
        RECT 949.265 172.405 975.920 172.415 ;
        RECT 1145.590 172.410 1172.245 172.420 ;
        RECT 537.825 172.130 556.730 172.140 ;
        RECT 734.190 172.135 753.095 172.145 ;
        RECT 930.575 172.130 975.920 172.405 ;
        RECT 1126.900 172.135 1172.245 172.410 ;
        RECT 930.575 172.120 949.480 172.130 ;
        RECT 1126.900 172.125 1145.805 172.135 ;
        RECT 341.505 172.085 360.410 172.095 ;
        RECT 188.450 170.970 188.830 171.005 ;
        RECT 581.160 170.975 581.540 171.010 ;
        RECT 777.525 170.980 777.905 171.015 ;
        RECT -58.045 170.880 -57.665 170.915 ;
        RECT -79.545 170.775 -79.165 170.815 ;
        RECT -79.615 170.470 -76.780 170.775 ;
        RECT -60.800 170.570 -57.665 170.880 ;
        RECT 166.950 170.865 167.330 170.905 ;
        RECT -58.045 170.535 -57.665 170.570 ;
        RECT 166.880 170.560 169.715 170.865 ;
        RECT 185.695 170.660 188.830 170.970 ;
        RECT 384.840 170.930 385.220 170.965 ;
        RECT 363.340 170.825 363.720 170.865 ;
        RECT 188.450 170.625 188.830 170.660 ;
        RECT 166.950 170.525 167.330 170.560 ;
        RECT 363.270 170.520 366.105 170.825 ;
        RECT 382.085 170.620 385.220 170.930 ;
        RECT 559.660 170.870 560.040 170.910 ;
        RECT 384.840 170.585 385.220 170.620 ;
        RECT 559.590 170.565 562.425 170.870 ;
        RECT 578.405 170.665 581.540 170.975 ;
        RECT 756.025 170.875 756.405 170.915 ;
        RECT 581.160 170.630 581.540 170.665 ;
        RECT 755.955 170.570 758.790 170.875 ;
        RECT 774.770 170.670 777.905 170.980 ;
        RECT 973.910 170.965 974.290 171.000 ;
        RECT 1170.235 170.970 1170.615 171.005 ;
        RECT 952.410 170.860 952.790 170.900 ;
        RECT 777.525 170.635 777.905 170.670 ;
        RECT 559.660 170.530 560.040 170.565 ;
        RECT 756.025 170.535 756.405 170.570 ;
        RECT 952.340 170.555 955.175 170.860 ;
        RECT 971.155 170.655 974.290 170.965 ;
        RECT 1148.735 170.865 1149.115 170.905 ;
        RECT 973.910 170.620 974.290 170.655 ;
        RECT 1148.665 170.560 1151.500 170.865 ;
        RECT 1167.480 170.660 1170.615 170.970 ;
        RECT 1170.235 170.625 1170.615 170.660 ;
        RECT 952.410 170.520 952.790 170.555 ;
        RECT 1148.735 170.525 1149.115 170.560 ;
        RECT 363.340 170.485 363.720 170.520 ;
        RECT -79.545 170.435 -79.165 170.470 ;
        RECT -75.545 162.645 -74.455 163.025 ;
        RECT -63.000 162.645 -61.665 163.025 ;
        RECT 170.950 162.735 172.040 163.115 ;
        RECT 183.495 162.735 184.830 163.115 ;
        RECT 367.340 162.695 368.430 163.075 ;
        RECT 379.885 162.695 381.220 163.075 ;
        RECT 563.660 162.740 564.750 163.120 ;
        RECT 576.205 162.740 577.540 163.120 ;
        RECT 760.025 162.745 761.115 163.125 ;
        RECT 772.570 162.745 773.905 163.125 ;
        RECT 956.410 162.730 957.500 163.110 ;
        RECT 968.955 162.730 970.290 163.110 ;
        RECT 1152.735 162.735 1153.825 163.115 ;
        RECT 1165.280 162.735 1166.615 163.115 ;
        RECT -75.060 160.650 -62.210 160.985 ;
        RECT 171.435 160.740 184.285 161.075 ;
        RECT 367.825 160.700 380.675 161.035 ;
        RECT 564.145 160.745 576.995 161.080 ;
        RECT 760.510 160.750 773.360 161.085 ;
        RECT 956.895 160.735 969.745 161.070 ;
        RECT 1153.220 160.740 1166.070 161.075 ;
      LAYER Metal2 ;
        RECT -100.700 18.030 -100.405 204.520 ;
        RECT -77.145 170.350 -76.855 172.410 ;
        RECT -74.855 160.435 -74.530 163.200 ;
        RECT -68.275 160.560 -67.985 172.395 ;
        RECT -60.370 170.290 -60.060 172.805 ;
        RECT -62.920 160.435 -62.595 163.200 ;
        RECT -50.940 17.775 -50.645 204.515 ;
        RECT -26.910 190.085 -26.620 192.145 ;
        RECT -24.620 180.170 -24.295 182.935 ;
        RECT -18.040 180.295 -17.750 192.130 ;
        RECT -10.135 190.025 -9.825 192.540 ;
        RECT -12.685 180.170 -12.360 182.935 ;
        RECT 145.230 17.785 145.525 204.525 ;
        RECT 169.350 170.440 169.640 172.500 ;
        RECT 171.640 160.525 171.965 163.290 ;
        RECT 178.220 160.650 178.510 172.485 ;
        RECT 186.125 170.380 186.435 172.895 ;
        RECT 183.575 160.525 183.900 163.290 ;
        RECT 341.620 17.745 341.915 204.485 ;
        RECT 365.740 170.400 366.030 172.460 ;
        RECT 368.030 160.485 368.355 163.250 ;
        RECT 374.610 160.610 374.900 172.445 ;
        RECT 382.515 170.340 382.825 172.855 ;
        RECT 379.965 160.485 380.290 163.250 ;
        RECT 537.940 17.790 538.235 204.530 ;
        RECT 562.060 170.445 562.350 172.505 ;
        RECT 564.350 160.530 564.675 163.295 ;
        RECT 570.930 160.655 571.220 172.490 ;
        RECT 578.835 170.385 579.145 172.900 ;
        RECT 576.285 160.530 576.610 163.295 ;
        RECT 734.305 17.795 734.600 204.535 ;
        RECT 758.425 170.450 758.715 172.510 ;
        RECT 760.715 160.535 761.040 163.300 ;
        RECT 767.295 160.660 767.585 172.495 ;
        RECT 775.200 170.390 775.510 172.905 ;
        RECT 772.650 160.535 772.975 163.300 ;
        RECT 930.690 17.780 930.985 204.520 ;
        RECT 954.810 170.435 955.100 172.495 ;
        RECT 957.100 160.520 957.425 163.285 ;
        RECT 963.680 160.645 963.970 172.480 ;
        RECT 971.585 170.375 971.895 172.890 ;
        RECT 969.035 160.520 969.360 163.285 ;
        RECT 1127.015 17.785 1127.310 204.525 ;
        RECT 1151.135 170.440 1151.425 172.500 ;
        RECT 1153.425 160.525 1153.750 163.290 ;
        RECT 1160.005 160.650 1160.295 172.485 ;
        RECT 1167.910 170.380 1168.220 172.895 ;
        RECT 1165.360 160.525 1165.685 163.290 ;
    END
  END b6_p0
  PIN b6_p1_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.575 201.445 1143.740 201.715 ;
        RECT -21.220 168.550 -20.840 168.595 ;
        RECT -15.720 168.550 -15.340 168.595 ;
        RECT -21.270 168.235 -15.335 168.550 ;
        RECT -21.220 168.215 -20.840 168.235 ;
        RECT -15.720 168.215 -15.340 168.235 ;
        RECT -29.220 160.725 -28.130 161.105 ;
        RECT -7.720 161.060 -7.340 161.105 ;
        RECT -8.455 160.760 -7.145 161.060 ;
        RECT -7.720 160.725 -7.340 160.760 ;
        RECT -48.120 160.215 -32.175 160.240 ;
        RECT -48.120 159.890 -5.710 160.215 ;
        RECT -32.365 159.865 -5.710 159.890 ;
        RECT 174.865 148.845 175.245 148.890 ;
        RECT 180.365 148.845 180.745 148.890 ;
        RECT 567.575 148.850 567.955 148.895 ;
        RECT 573.075 148.850 573.455 148.895 ;
        RECT 763.940 148.855 764.320 148.900 ;
        RECT 769.440 148.855 769.820 148.900 ;
        RECT -71.630 148.755 -71.250 148.800 ;
        RECT -66.130 148.755 -65.750 148.800 ;
        RECT -71.680 148.440 -65.745 148.755 ;
        RECT 174.815 148.530 180.750 148.845 ;
        RECT 371.255 148.805 371.635 148.850 ;
        RECT 376.755 148.805 377.135 148.850 ;
        RECT 174.865 148.510 175.245 148.530 ;
        RECT 180.365 148.510 180.745 148.530 ;
        RECT 371.205 148.490 377.140 148.805 ;
        RECT 567.525 148.535 573.460 148.850 ;
        RECT 763.890 148.540 769.825 148.855 ;
        RECT 960.325 148.840 960.705 148.885 ;
        RECT 965.825 148.840 966.205 148.885 ;
        RECT 1156.650 148.845 1157.030 148.890 ;
        RECT 1162.150 148.845 1162.530 148.890 ;
        RECT 567.575 148.515 567.955 148.535 ;
        RECT 573.075 148.515 573.455 148.535 ;
        RECT 763.940 148.520 764.320 148.540 ;
        RECT 769.440 148.520 769.820 148.540 ;
        RECT 960.275 148.525 966.210 148.840 ;
        RECT 1156.600 148.530 1162.535 148.845 ;
        RECT 960.325 148.505 960.705 148.525 ;
        RECT 965.825 148.505 966.205 148.525 ;
        RECT 1156.650 148.510 1157.030 148.530 ;
        RECT 1162.150 148.510 1162.530 148.530 ;
        RECT 371.255 148.470 371.635 148.490 ;
        RECT 376.755 148.470 377.135 148.490 ;
        RECT -71.630 148.420 -71.250 148.440 ;
        RECT -66.130 148.420 -65.750 148.440 ;
        RECT -79.630 140.930 -78.540 141.310 ;
        RECT -58.130 141.265 -57.750 141.310 ;
        RECT -58.865 140.965 -57.555 141.265 ;
        RECT 166.865 141.020 167.955 141.400 ;
        RECT 188.365 141.355 188.745 141.400 ;
        RECT 187.630 141.055 188.940 141.355 ;
        RECT 188.365 141.020 188.745 141.055 ;
        RECT 363.255 140.980 364.345 141.360 ;
        RECT 384.755 141.315 385.135 141.360 ;
        RECT 384.020 141.015 385.330 141.315 ;
        RECT 559.575 141.025 560.665 141.405 ;
        RECT 581.075 141.360 581.455 141.405 ;
        RECT 580.340 141.060 581.650 141.360 ;
        RECT 581.075 141.025 581.455 141.060 ;
        RECT 755.940 141.030 757.030 141.410 ;
        RECT 777.440 141.365 777.820 141.410 ;
        RECT 776.705 141.065 778.015 141.365 ;
        RECT 777.440 141.030 777.820 141.065 ;
        RECT 952.325 141.015 953.415 141.395 ;
        RECT 973.825 141.350 974.205 141.395 ;
        RECT 973.090 141.050 974.400 141.350 ;
        RECT 973.825 141.015 974.205 141.050 ;
        RECT 1148.650 141.020 1149.740 141.400 ;
        RECT 1170.150 141.355 1170.530 141.400 ;
        RECT 1169.415 141.055 1170.725 141.355 ;
        RECT 1170.150 141.020 1170.530 141.055 ;
        RECT 384.755 140.980 385.135 141.015 ;
        RECT -58.130 140.930 -57.750 140.965 ;
        RECT 148.040 140.510 163.985 140.520 ;
        RECT 540.750 140.515 556.695 140.525 ;
        RECT 737.115 140.520 753.060 140.530 ;
        RECT -97.885 140.070 -56.120 140.420 ;
        RECT 148.040 140.170 190.375 140.510 ;
        RECT 163.720 140.160 190.375 140.170 ;
        RECT 344.430 140.470 360.375 140.480 ;
        RECT 344.430 140.130 386.765 140.470 ;
        RECT 540.750 140.175 583.085 140.515 ;
        RECT 737.115 140.180 779.450 140.520 ;
        RECT 556.430 140.165 583.085 140.175 ;
        RECT 752.795 140.170 779.450 140.180 ;
        RECT 933.500 140.505 949.445 140.515 ;
        RECT 1129.825 140.510 1145.770 140.520 ;
        RECT 933.500 140.165 975.835 140.505 ;
        RECT 1129.825 140.170 1172.160 140.510 ;
        RECT 949.180 140.155 975.835 140.165 ;
        RECT 1145.505 140.160 1172.160 140.170 ;
        RECT 360.110 140.120 386.765 140.130 ;
      LAYER Metal2 ;
        RECT -97.710 18.040 -97.420 204.530 ;
        RECT -79.015 140.070 -78.635 141.445 ;
        RECT -69.305 139.780 -68.935 148.880 ;
        RECT -58.760 139.985 -58.425 141.335 ;
        RECT -47.950 17.885 -47.660 204.500 ;
        RECT -28.605 159.865 -28.225 161.240 ;
        RECT -18.895 159.575 -18.525 168.675 ;
        RECT -8.350 159.780 -8.015 161.130 ;
        RECT 148.220 17.895 148.510 204.510 ;
        RECT 167.480 140.160 167.860 141.535 ;
        RECT 177.190 139.870 177.560 148.970 ;
        RECT 187.735 140.075 188.070 141.425 ;
        RECT 344.610 17.855 344.900 204.470 ;
        RECT 363.870 140.120 364.250 141.495 ;
        RECT 373.580 139.830 373.950 148.930 ;
        RECT 384.125 140.035 384.460 141.385 ;
        RECT 540.930 17.900 541.220 204.515 ;
        RECT 560.190 140.165 560.570 141.540 ;
        RECT 569.900 139.875 570.270 148.975 ;
        RECT 580.445 140.080 580.780 141.430 ;
        RECT 737.295 17.905 737.585 204.520 ;
        RECT 756.555 140.170 756.935 141.545 ;
        RECT 766.265 139.880 766.635 148.980 ;
        RECT 776.810 140.085 777.145 141.435 ;
        RECT 933.680 17.890 933.970 204.505 ;
        RECT 952.940 140.155 953.320 141.530 ;
        RECT 962.650 139.865 963.020 148.965 ;
        RECT 973.195 140.070 973.530 141.420 ;
        RECT 1130.005 17.895 1130.295 204.510 ;
        RECT 1149.265 140.160 1149.645 141.535 ;
        RECT 1158.975 139.870 1159.345 148.970 ;
        RECT 1169.520 140.075 1169.855 141.425 ;
    END
  END b6_p1_not
  PIN b6_p1
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.605 201.965 1143.740 202.255 ;
        RECT -49.090 172.410 -32.175 172.435 ;
        RECT -49.090 172.150 -5.710 172.410 ;
        RECT -32.365 172.125 -5.710 172.150 ;
        RECT -7.720 170.960 -7.340 170.995 ;
        RECT -29.220 170.855 -28.840 170.895 ;
        RECT -29.290 170.550 -26.455 170.855 ;
        RECT -10.475 170.650 -7.340 170.960 ;
        RECT -7.720 170.615 -7.340 170.650 ;
        RECT -29.220 170.515 -28.840 170.550 ;
        RECT -25.220 162.725 -24.130 163.105 ;
        RECT -12.675 162.725 -11.340 163.105 ;
        RECT -24.735 160.730 -11.885 161.065 ;
        RECT 147.070 152.705 163.985 152.715 ;
        RECT 539.780 152.710 556.695 152.720 ;
        RECT 736.145 152.715 753.060 152.725 ;
        RECT -98.855 152.330 -56.120 152.615 ;
        RECT 147.070 152.430 190.375 152.705 ;
        RECT 163.720 152.420 190.375 152.430 ;
        RECT 343.460 152.665 360.375 152.675 ;
        RECT 343.460 152.390 386.765 152.665 ;
        RECT 539.780 152.435 583.085 152.710 ;
        RECT 736.145 152.440 779.450 152.715 ;
        RECT 556.430 152.425 583.085 152.435 ;
        RECT 752.795 152.430 779.450 152.440 ;
        RECT 932.530 152.700 949.445 152.710 ;
        RECT 1128.855 152.705 1145.770 152.715 ;
        RECT 932.530 152.425 975.835 152.700 ;
        RECT 1128.855 152.430 1172.160 152.705 ;
        RECT 949.180 152.415 975.835 152.425 ;
        RECT 1145.505 152.420 1172.160 152.430 ;
        RECT 360.110 152.380 386.765 152.390 ;
        RECT 188.365 151.255 188.745 151.290 ;
        RECT 581.075 151.260 581.455 151.295 ;
        RECT 777.440 151.265 777.820 151.300 ;
        RECT -58.130 151.165 -57.750 151.200 ;
        RECT -79.630 151.060 -79.250 151.100 ;
        RECT -79.700 150.755 -76.865 151.060 ;
        RECT -60.885 150.855 -57.750 151.165 ;
        RECT 166.865 151.150 167.245 151.190 ;
        RECT -58.130 150.820 -57.750 150.855 ;
        RECT 166.795 150.845 169.630 151.150 ;
        RECT 185.610 150.945 188.745 151.255 ;
        RECT 384.755 151.215 385.135 151.250 ;
        RECT 363.255 151.110 363.635 151.150 ;
        RECT 188.365 150.910 188.745 150.945 ;
        RECT 166.865 150.810 167.245 150.845 ;
        RECT 363.185 150.805 366.020 151.110 ;
        RECT 382.000 150.905 385.135 151.215 ;
        RECT 559.575 151.155 559.955 151.195 ;
        RECT 384.755 150.870 385.135 150.905 ;
        RECT 559.505 150.850 562.340 151.155 ;
        RECT 578.320 150.950 581.455 151.260 ;
        RECT 755.940 151.160 756.320 151.200 ;
        RECT 581.075 150.915 581.455 150.950 ;
        RECT 755.870 150.855 758.705 151.160 ;
        RECT 774.685 150.955 777.820 151.265 ;
        RECT 973.825 151.250 974.205 151.285 ;
        RECT 1170.150 151.255 1170.530 151.290 ;
        RECT 952.325 151.145 952.705 151.185 ;
        RECT 777.440 150.920 777.820 150.955 ;
        RECT 559.575 150.815 559.955 150.850 ;
        RECT 755.940 150.820 756.320 150.855 ;
        RECT 952.255 150.840 955.090 151.145 ;
        RECT 971.070 150.940 974.205 151.250 ;
        RECT 1148.650 151.150 1149.030 151.190 ;
        RECT 973.825 150.905 974.205 150.940 ;
        RECT 1148.580 150.845 1151.415 151.150 ;
        RECT 1167.395 150.945 1170.530 151.255 ;
        RECT 1170.150 150.910 1170.530 150.945 ;
        RECT 952.325 150.805 952.705 150.840 ;
        RECT 1148.650 150.810 1149.030 150.845 ;
        RECT 363.255 150.770 363.635 150.805 ;
        RECT -79.630 150.720 -79.250 150.755 ;
        RECT -75.630 142.930 -74.540 143.310 ;
        RECT -63.085 142.930 -61.750 143.310 ;
        RECT 170.865 143.020 171.955 143.400 ;
        RECT 183.410 143.020 184.745 143.400 ;
        RECT 367.255 142.980 368.345 143.360 ;
        RECT 379.800 142.980 381.135 143.360 ;
        RECT 563.575 143.025 564.665 143.405 ;
        RECT 576.120 143.025 577.455 143.405 ;
        RECT 759.940 143.030 761.030 143.410 ;
        RECT 772.485 143.030 773.820 143.410 ;
        RECT 956.325 143.015 957.415 143.395 ;
        RECT 968.870 143.015 970.205 143.395 ;
        RECT 1152.650 143.020 1153.740 143.400 ;
        RECT 1165.195 143.020 1166.530 143.400 ;
        RECT -75.145 140.935 -62.295 141.270 ;
        RECT 171.350 141.025 184.200 141.360 ;
        RECT 367.740 140.985 380.590 141.320 ;
        RECT 564.060 141.030 576.910 141.365 ;
        RECT 760.425 141.035 773.275 141.370 ;
        RECT 956.810 141.020 969.660 141.355 ;
        RECT 1153.135 141.025 1165.985 141.360 ;
      LAYER Metal2 ;
        RECT -98.705 18.045 -98.415 204.525 ;
        RECT -77.230 150.635 -76.940 152.695 ;
        RECT -74.940 140.720 -74.615 143.485 ;
        RECT -68.360 140.845 -68.070 152.680 ;
        RECT -60.455 150.575 -60.145 153.090 ;
        RECT -63.005 140.720 -62.680 143.485 ;
        RECT -48.945 17.945 -48.655 204.515 ;
        RECT -26.820 170.430 -26.530 172.490 ;
        RECT -24.530 160.515 -24.205 163.280 ;
        RECT -17.950 160.640 -17.660 172.475 ;
        RECT -10.045 170.370 -9.735 172.885 ;
        RECT -12.595 160.515 -12.270 163.280 ;
        RECT 147.225 17.955 147.515 204.525 ;
        RECT 169.265 150.725 169.555 152.785 ;
        RECT 171.555 140.810 171.880 143.575 ;
        RECT 178.135 140.935 178.425 152.770 ;
        RECT 186.040 150.665 186.350 153.180 ;
        RECT 183.490 140.810 183.815 143.575 ;
        RECT 343.615 17.915 343.905 204.485 ;
        RECT 365.655 150.685 365.945 152.745 ;
        RECT 367.945 140.770 368.270 143.535 ;
        RECT 374.525 140.895 374.815 152.730 ;
        RECT 382.430 150.625 382.740 153.140 ;
        RECT 379.880 140.770 380.205 143.535 ;
        RECT 539.935 17.960 540.225 204.530 ;
        RECT 561.975 150.730 562.265 152.790 ;
        RECT 564.265 140.815 564.590 143.580 ;
        RECT 570.845 140.940 571.135 152.775 ;
        RECT 578.750 150.670 579.060 153.185 ;
        RECT 576.200 140.815 576.525 143.580 ;
        RECT 736.300 17.965 736.590 204.535 ;
        RECT 758.340 150.735 758.630 152.795 ;
        RECT 760.630 140.820 760.955 143.585 ;
        RECT 767.210 140.945 767.500 152.780 ;
        RECT 775.115 150.675 775.425 153.190 ;
        RECT 772.565 140.820 772.890 143.585 ;
        RECT 932.685 17.950 932.975 204.520 ;
        RECT 954.725 150.720 955.015 152.780 ;
        RECT 957.015 140.805 957.340 143.570 ;
        RECT 963.595 140.930 963.885 152.765 ;
        RECT 971.500 150.660 971.810 153.175 ;
        RECT 968.950 140.805 969.275 143.570 ;
        RECT 1129.010 17.955 1129.300 204.525 ;
        RECT 1151.050 150.725 1151.340 152.785 ;
        RECT 1153.340 140.810 1153.665 143.575 ;
        RECT 1159.920 140.935 1160.210 152.770 ;
        RECT 1167.825 150.665 1168.135 153.180 ;
        RECT 1165.275 140.810 1165.600 143.575 ;
    END
  END b6_p1
  PIN b6_p2_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.585 200.250 1143.745 200.575 ;
        RECT -21.305 148.835 -20.925 148.880 ;
        RECT -15.805 148.835 -15.425 148.880 ;
        RECT -21.355 148.520 -15.420 148.835 ;
        RECT -21.305 148.500 -20.925 148.520 ;
        RECT -15.805 148.500 -15.425 148.520 ;
        RECT -29.305 141.010 -28.215 141.390 ;
        RECT -7.805 141.345 -7.425 141.390 ;
        RECT -8.540 141.045 -7.230 141.345 ;
        RECT -7.805 141.010 -7.425 141.045 ;
        RECT -32.450 140.430 -5.795 140.500 ;
        RECT -46.080 140.150 -5.795 140.430 ;
        RECT -46.080 140.080 -32.005 140.150 ;
        RECT 174.925 129.040 175.305 129.085 ;
        RECT 180.425 129.040 180.805 129.085 ;
        RECT 567.635 129.045 568.015 129.090 ;
        RECT 573.135 129.045 573.515 129.090 ;
        RECT 764.000 129.050 764.380 129.095 ;
        RECT 769.500 129.050 769.880 129.095 ;
        RECT -71.570 128.950 -71.190 128.995 ;
        RECT -66.070 128.950 -65.690 128.995 ;
        RECT -71.620 128.635 -65.685 128.950 ;
        RECT 174.875 128.725 180.810 129.040 ;
        RECT 371.315 129.000 371.695 129.045 ;
        RECT 376.815 129.000 377.195 129.045 ;
        RECT 174.925 128.705 175.305 128.725 ;
        RECT 180.425 128.705 180.805 128.725 ;
        RECT 371.265 128.685 377.200 129.000 ;
        RECT 567.585 128.730 573.520 129.045 ;
        RECT 763.950 128.735 769.885 129.050 ;
        RECT 960.385 129.035 960.765 129.080 ;
        RECT 965.885 129.035 966.265 129.080 ;
        RECT 1156.710 129.040 1157.090 129.085 ;
        RECT 1162.210 129.040 1162.590 129.085 ;
        RECT 567.635 128.710 568.015 128.730 ;
        RECT 573.135 128.710 573.515 128.730 ;
        RECT 764.000 128.715 764.380 128.735 ;
        RECT 769.500 128.715 769.880 128.735 ;
        RECT 960.335 128.720 966.270 129.035 ;
        RECT 1156.660 128.725 1162.595 129.040 ;
        RECT 960.385 128.700 960.765 128.720 ;
        RECT 965.885 128.700 966.265 128.720 ;
        RECT 1156.710 128.705 1157.090 128.725 ;
        RECT 1162.210 128.705 1162.590 128.725 ;
        RECT 371.315 128.665 371.695 128.685 ;
        RECT 376.815 128.665 377.195 128.685 ;
        RECT -71.570 128.615 -71.190 128.635 ;
        RECT -66.070 128.615 -65.690 128.635 ;
        RECT -79.570 121.125 -78.480 121.505 ;
        RECT -58.070 121.460 -57.690 121.505 ;
        RECT -58.805 121.160 -57.495 121.460 ;
        RECT 166.925 121.215 168.015 121.595 ;
        RECT 188.425 121.550 188.805 121.595 ;
        RECT 187.690 121.250 189.000 121.550 ;
        RECT 188.425 121.215 188.805 121.250 ;
        RECT 363.315 121.175 364.405 121.555 ;
        RECT 384.815 121.510 385.195 121.555 ;
        RECT 384.080 121.210 385.390 121.510 ;
        RECT 559.635 121.220 560.725 121.600 ;
        RECT 581.135 121.555 581.515 121.600 ;
        RECT 580.400 121.255 581.710 121.555 ;
        RECT 581.135 121.220 581.515 121.255 ;
        RECT 756.000 121.225 757.090 121.605 ;
        RECT 777.500 121.560 777.880 121.605 ;
        RECT 776.765 121.260 778.075 121.560 ;
        RECT 777.500 121.225 777.880 121.260 ;
        RECT 952.385 121.210 953.475 121.590 ;
        RECT 973.885 121.545 974.265 121.590 ;
        RECT 973.150 121.245 974.460 121.545 ;
        RECT 973.885 121.210 974.265 121.245 ;
        RECT 1148.710 121.215 1149.800 121.595 ;
        RECT 1170.210 121.550 1170.590 121.595 ;
        RECT 1169.475 121.250 1170.785 121.550 ;
        RECT 1170.210 121.215 1170.590 121.250 ;
        RECT 384.815 121.175 385.195 121.210 ;
        RECT -58.070 121.125 -57.690 121.160 ;
        RECT 739.155 120.715 753.230 120.720 ;
        RECT 542.790 120.710 556.865 120.715 ;
        RECT 150.080 120.705 164.155 120.710 ;
        RECT -82.715 120.610 -56.060 120.615 ;
        RECT -95.845 120.265 -56.060 120.610 ;
        RECT 150.080 120.360 190.435 120.705 ;
        RECT 163.780 120.355 190.435 120.360 ;
        RECT 346.470 120.665 360.545 120.670 ;
        RECT 346.470 120.320 386.825 120.665 ;
        RECT 542.790 120.365 583.145 120.710 ;
        RECT 739.155 120.370 779.510 120.715 ;
        RECT 1131.865 120.705 1145.940 120.710 ;
        RECT 752.855 120.365 779.510 120.370 ;
        RECT 935.540 120.700 949.615 120.705 ;
        RECT 556.490 120.360 583.145 120.365 ;
        RECT 935.540 120.355 975.895 120.700 ;
        RECT 1131.865 120.360 1172.220 120.705 ;
        RECT 1145.565 120.355 1172.220 120.360 ;
        RECT 949.240 120.350 975.895 120.355 ;
        RECT 360.170 120.315 386.825 120.320 ;
        RECT -95.845 120.260 -82.555 120.265 ;
      LAYER Metal2 ;
        RECT -95.655 18.040 -95.205 204.535 ;
        RECT -78.955 120.265 -78.575 121.640 ;
        RECT -69.245 119.975 -68.875 129.075 ;
        RECT -58.700 120.180 -58.365 121.530 ;
        RECT -45.895 18.025 -45.445 204.500 ;
        RECT -28.690 140.150 -28.310 141.525 ;
        RECT -18.980 139.860 -18.610 148.960 ;
        RECT -8.435 140.065 -8.100 141.415 ;
        RECT 150.275 18.035 150.725 204.510 ;
        RECT 167.540 120.355 167.920 121.730 ;
        RECT 177.250 120.065 177.620 129.165 ;
        RECT 187.795 120.270 188.130 121.620 ;
        RECT 346.665 17.995 347.115 204.470 ;
        RECT 363.930 120.315 364.310 121.690 ;
        RECT 373.640 120.025 374.010 129.125 ;
        RECT 384.185 120.230 384.520 121.580 ;
        RECT 542.985 18.040 543.435 204.515 ;
        RECT 560.250 120.360 560.630 121.735 ;
        RECT 569.960 120.070 570.330 129.170 ;
        RECT 580.505 120.275 580.840 121.625 ;
        RECT 739.350 18.045 739.800 204.520 ;
        RECT 756.615 120.365 756.995 121.740 ;
        RECT 766.325 120.075 766.695 129.175 ;
        RECT 776.870 120.280 777.205 121.630 ;
        RECT 935.735 18.030 936.185 204.505 ;
        RECT 953.000 120.350 953.380 121.725 ;
        RECT 962.710 120.060 963.080 129.160 ;
        RECT 973.255 120.265 973.590 121.615 ;
        RECT 1132.060 18.035 1132.510 204.510 ;
        RECT 1149.325 120.355 1149.705 121.730 ;
        RECT 1159.035 120.065 1159.405 129.165 ;
        RECT 1169.580 120.270 1169.915 121.620 ;
    END
  END b6_p2_not
  PIN b6_p2
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.560 200.885 1143.755 201.160 ;
        RECT -32.450 152.625 -5.795 152.695 ;
        RECT -47.145 152.410 -5.795 152.625 ;
        RECT -47.145 152.340 -31.975 152.410 ;
        RECT -7.805 151.245 -7.425 151.280 ;
        RECT -29.305 151.140 -28.925 151.180 ;
        RECT -29.375 150.835 -26.540 151.140 ;
        RECT -10.560 150.935 -7.425 151.245 ;
        RECT -7.805 150.900 -7.425 150.935 ;
        RECT -29.305 150.800 -28.925 150.835 ;
        RECT -25.305 143.010 -24.215 143.390 ;
        RECT -12.760 143.010 -11.425 143.390 ;
        RECT -24.820 141.015 -11.970 141.350 ;
        RECT 738.090 132.910 753.260 132.915 ;
        RECT 541.725 132.905 556.895 132.910 ;
        RECT 149.015 132.900 164.185 132.905 ;
        RECT -82.715 132.805 -56.060 132.810 ;
        RECT -96.910 132.525 -56.060 132.805 ;
        RECT 149.015 132.620 190.435 132.900 ;
        RECT 163.780 132.615 190.435 132.620 ;
        RECT 345.405 132.860 360.575 132.865 ;
        RECT 345.405 132.580 386.825 132.860 ;
        RECT 541.725 132.625 583.145 132.905 ;
        RECT 738.090 132.630 779.510 132.910 ;
        RECT 1130.800 132.900 1145.970 132.905 ;
        RECT 752.855 132.625 779.510 132.630 ;
        RECT 934.475 132.895 949.645 132.900 ;
        RECT 556.490 132.620 583.145 132.625 ;
        RECT 934.475 132.615 975.895 132.895 ;
        RECT 1130.800 132.620 1172.220 132.900 ;
        RECT 1145.565 132.615 1172.220 132.620 ;
        RECT 949.240 132.610 975.895 132.615 ;
        RECT 360.170 132.575 386.825 132.580 ;
        RECT -96.910 132.520 -82.455 132.525 ;
        RECT 188.425 131.450 188.805 131.485 ;
        RECT 581.135 131.455 581.515 131.490 ;
        RECT 777.500 131.460 777.880 131.495 ;
        RECT -58.070 131.360 -57.690 131.395 ;
        RECT -79.570 131.255 -79.190 131.295 ;
        RECT -79.640 130.950 -76.805 131.255 ;
        RECT -60.825 131.050 -57.690 131.360 ;
        RECT 166.925 131.345 167.305 131.385 ;
        RECT -58.070 131.015 -57.690 131.050 ;
        RECT 166.855 131.040 169.690 131.345 ;
        RECT 185.670 131.140 188.805 131.450 ;
        RECT 384.815 131.410 385.195 131.445 ;
        RECT 363.315 131.305 363.695 131.345 ;
        RECT 188.425 131.105 188.805 131.140 ;
        RECT 166.925 131.005 167.305 131.040 ;
        RECT 363.245 131.000 366.080 131.305 ;
        RECT 382.060 131.100 385.195 131.410 ;
        RECT 559.635 131.350 560.015 131.390 ;
        RECT 384.815 131.065 385.195 131.100 ;
        RECT 559.565 131.045 562.400 131.350 ;
        RECT 578.380 131.145 581.515 131.455 ;
        RECT 756.000 131.355 756.380 131.395 ;
        RECT 581.135 131.110 581.515 131.145 ;
        RECT 755.930 131.050 758.765 131.355 ;
        RECT 774.745 131.150 777.880 131.460 ;
        RECT 973.885 131.445 974.265 131.480 ;
        RECT 1170.210 131.450 1170.590 131.485 ;
        RECT 952.385 131.340 952.765 131.380 ;
        RECT 777.500 131.115 777.880 131.150 ;
        RECT 559.635 131.010 560.015 131.045 ;
        RECT 756.000 131.015 756.380 131.050 ;
        RECT 952.315 131.035 955.150 131.340 ;
        RECT 971.130 131.135 974.265 131.445 ;
        RECT 1148.710 131.345 1149.090 131.385 ;
        RECT 973.885 131.100 974.265 131.135 ;
        RECT 1148.640 131.040 1151.475 131.345 ;
        RECT 1167.455 131.140 1170.590 131.450 ;
        RECT 1170.210 131.105 1170.590 131.140 ;
        RECT 952.385 131.000 952.765 131.035 ;
        RECT 1148.710 131.005 1149.090 131.040 ;
        RECT 363.315 130.965 363.695 131.000 ;
        RECT -79.570 130.915 -79.190 130.950 ;
        RECT -75.570 123.125 -74.480 123.505 ;
        RECT -63.025 123.125 -61.690 123.505 ;
        RECT 170.925 123.215 172.015 123.595 ;
        RECT 183.470 123.215 184.805 123.595 ;
        RECT 367.315 123.175 368.405 123.555 ;
        RECT 379.860 123.175 381.195 123.555 ;
        RECT 563.635 123.220 564.725 123.600 ;
        RECT 576.180 123.220 577.515 123.600 ;
        RECT 760.000 123.225 761.090 123.605 ;
        RECT 772.545 123.225 773.880 123.605 ;
        RECT 956.385 123.210 957.475 123.590 ;
        RECT 968.930 123.210 970.265 123.590 ;
        RECT 1152.710 123.215 1153.800 123.595 ;
        RECT 1165.255 123.215 1166.590 123.595 ;
        RECT -75.085 121.130 -62.235 121.465 ;
        RECT 171.410 121.220 184.260 121.555 ;
        RECT 367.800 121.180 380.650 121.515 ;
        RECT 564.120 121.225 576.970 121.560 ;
        RECT 760.485 121.230 773.335 121.565 ;
        RECT 956.870 121.215 969.720 121.550 ;
        RECT 1153.195 121.220 1166.045 121.555 ;
      LAYER Metal2 ;
        RECT -96.750 18.040 -96.425 204.535 ;
        RECT -77.170 130.830 -76.880 132.890 ;
        RECT -74.880 120.915 -74.555 123.680 ;
        RECT -68.300 121.040 -68.010 132.875 ;
        RECT -60.395 130.770 -60.085 133.285 ;
        RECT -62.945 120.915 -62.620 123.680 ;
        RECT -46.990 17.990 -46.665 204.515 ;
        RECT -26.905 150.715 -26.615 152.775 ;
        RECT -24.615 140.800 -24.290 143.565 ;
        RECT -18.035 140.925 -17.745 152.760 ;
        RECT -10.130 150.655 -9.820 153.170 ;
        RECT -12.680 140.800 -12.355 143.565 ;
        RECT 149.180 18.000 149.505 204.525 ;
        RECT 169.325 130.920 169.615 132.980 ;
        RECT 171.615 121.005 171.940 123.770 ;
        RECT 178.195 121.130 178.485 132.965 ;
        RECT 186.100 130.860 186.410 133.375 ;
        RECT 183.550 121.005 183.875 123.770 ;
        RECT 345.570 17.960 345.895 204.485 ;
        RECT 365.715 130.880 366.005 132.940 ;
        RECT 368.005 120.965 368.330 123.730 ;
        RECT 374.585 121.090 374.875 132.925 ;
        RECT 382.490 130.820 382.800 133.335 ;
        RECT 379.940 120.965 380.265 123.730 ;
        RECT 541.890 18.005 542.215 204.530 ;
        RECT 562.035 130.925 562.325 132.985 ;
        RECT 564.325 121.010 564.650 123.775 ;
        RECT 570.905 121.135 571.195 132.970 ;
        RECT 578.810 130.865 579.120 133.380 ;
        RECT 576.260 121.010 576.585 123.775 ;
        RECT 738.255 18.010 738.580 204.535 ;
        RECT 758.400 130.930 758.690 132.990 ;
        RECT 760.690 121.015 761.015 123.780 ;
        RECT 767.270 121.140 767.560 132.975 ;
        RECT 775.175 130.870 775.485 133.385 ;
        RECT 772.625 121.015 772.950 123.780 ;
        RECT 934.640 17.995 934.965 204.520 ;
        RECT 954.785 130.915 955.075 132.975 ;
        RECT 957.075 121.000 957.400 123.765 ;
        RECT 963.655 121.125 963.945 132.960 ;
        RECT 971.560 130.855 971.870 133.370 ;
        RECT 969.010 121.000 969.335 123.765 ;
        RECT 1130.965 18.000 1131.290 204.525 ;
        RECT 1151.110 130.920 1151.400 132.980 ;
        RECT 1153.400 121.005 1153.725 123.770 ;
        RECT 1159.980 121.130 1160.270 132.965 ;
        RECT 1167.885 130.860 1168.195 133.375 ;
        RECT 1165.335 121.005 1165.660 123.770 ;
    END
  END b6_p2
  PIN b6_p3
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.655 199.595 1143.755 199.910 ;
        RECT -32.390 132.865 -5.735 132.890 ;
        RECT -44.760 132.605 -5.735 132.865 ;
        RECT -44.760 132.580 -32.235 132.605 ;
        RECT -7.745 131.440 -7.365 131.475 ;
        RECT -29.245 131.335 -28.865 131.375 ;
        RECT -29.315 131.030 -26.480 131.335 ;
        RECT -10.500 131.130 -7.365 131.440 ;
        RECT -7.745 131.095 -7.365 131.130 ;
        RECT -29.245 130.995 -28.865 131.030 ;
        RECT -25.245 123.205 -24.155 123.585 ;
        RECT -12.700 123.205 -11.365 123.585 ;
        RECT -24.760 121.210 -11.910 121.545 ;
        RECT 151.400 113.130 163.925 113.145 ;
        RECT 544.110 113.135 556.635 113.150 ;
        RECT 740.475 113.140 753.000 113.155 ;
        RECT -94.525 113.040 -82.450 113.045 ;
        RECT -94.525 112.760 -56.130 113.040 ;
        RECT 151.400 112.860 190.365 113.130 ;
        RECT 163.710 112.845 190.365 112.860 ;
        RECT 347.790 113.090 360.315 113.105 ;
        RECT 347.790 112.820 386.755 113.090 ;
        RECT 544.110 112.865 583.075 113.135 ;
        RECT 740.475 112.870 779.440 113.140 ;
        RECT 556.420 112.850 583.075 112.865 ;
        RECT 752.785 112.855 779.440 112.870 ;
        RECT 936.860 113.125 949.385 113.140 ;
        RECT 1133.185 113.130 1145.710 113.145 ;
        RECT 936.860 112.855 975.825 113.125 ;
        RECT 1133.185 112.860 1172.150 113.130 ;
        RECT 949.170 112.840 975.825 112.855 ;
        RECT 1145.495 112.845 1172.150 112.860 ;
        RECT 360.100 112.805 386.755 112.820 ;
        RECT -82.785 112.755 -56.130 112.760 ;
        RECT 188.355 111.680 188.735 111.715 ;
        RECT 581.065 111.685 581.445 111.720 ;
        RECT 777.430 111.690 777.810 111.725 ;
        RECT -58.140 111.590 -57.760 111.625 ;
        RECT -79.640 111.485 -79.260 111.525 ;
        RECT -79.710 111.180 -76.875 111.485 ;
        RECT -60.895 111.280 -57.760 111.590 ;
        RECT 166.855 111.575 167.235 111.615 ;
        RECT -58.140 111.245 -57.760 111.280 ;
        RECT 166.785 111.270 169.620 111.575 ;
        RECT 185.600 111.370 188.735 111.680 ;
        RECT 384.745 111.640 385.125 111.675 ;
        RECT 363.245 111.535 363.625 111.575 ;
        RECT 188.355 111.335 188.735 111.370 ;
        RECT 166.855 111.235 167.235 111.270 ;
        RECT 363.175 111.230 366.010 111.535 ;
        RECT 381.990 111.330 385.125 111.640 ;
        RECT 559.565 111.580 559.945 111.620 ;
        RECT 384.745 111.295 385.125 111.330 ;
        RECT 559.495 111.275 562.330 111.580 ;
        RECT 578.310 111.375 581.445 111.685 ;
        RECT 755.930 111.585 756.310 111.625 ;
        RECT 581.065 111.340 581.445 111.375 ;
        RECT 755.860 111.280 758.695 111.585 ;
        RECT 774.675 111.380 777.810 111.690 ;
        RECT 973.815 111.675 974.195 111.710 ;
        RECT 1170.140 111.680 1170.520 111.715 ;
        RECT 952.315 111.570 952.695 111.610 ;
        RECT 777.430 111.345 777.810 111.380 ;
        RECT 559.565 111.240 559.945 111.275 ;
        RECT 755.930 111.245 756.310 111.280 ;
        RECT 952.245 111.265 955.080 111.570 ;
        RECT 971.060 111.365 974.195 111.675 ;
        RECT 1148.640 111.575 1149.020 111.615 ;
        RECT 973.815 111.330 974.195 111.365 ;
        RECT 1148.570 111.270 1151.405 111.575 ;
        RECT 1167.385 111.370 1170.520 111.680 ;
        RECT 1170.140 111.335 1170.520 111.370 ;
        RECT 952.315 111.230 952.695 111.265 ;
        RECT 1148.640 111.235 1149.020 111.270 ;
        RECT 363.245 111.195 363.625 111.230 ;
        RECT -79.640 111.145 -79.260 111.180 ;
        RECT -75.640 103.355 -74.550 103.735 ;
        RECT -63.095 103.355 -61.760 103.735 ;
        RECT 170.855 103.445 171.945 103.825 ;
        RECT 183.400 103.445 184.735 103.825 ;
        RECT 367.245 103.405 368.335 103.785 ;
        RECT 379.790 103.405 381.125 103.785 ;
        RECT 563.565 103.450 564.655 103.830 ;
        RECT 576.110 103.450 577.445 103.830 ;
        RECT 759.930 103.455 761.020 103.835 ;
        RECT 772.475 103.455 773.810 103.835 ;
        RECT 956.315 103.440 957.405 103.820 ;
        RECT 968.860 103.440 970.195 103.820 ;
        RECT 1152.640 103.445 1153.730 103.825 ;
        RECT 1165.185 103.445 1166.520 103.825 ;
        RECT -75.155 101.360 -62.305 101.695 ;
        RECT 171.340 101.450 184.190 101.785 ;
        RECT 367.730 101.410 380.580 101.745 ;
        RECT 564.050 101.455 576.900 101.790 ;
        RECT 760.415 101.460 773.265 101.795 ;
        RECT 956.800 101.445 969.650 101.780 ;
        RECT 1153.125 101.450 1165.975 101.785 ;
      LAYER Metal2 ;
        RECT -94.370 18.040 -94.010 204.520 ;
        RECT -77.240 111.060 -76.950 113.120 ;
        RECT -74.950 101.145 -74.625 103.910 ;
        RECT -68.370 101.270 -68.080 113.105 ;
        RECT -60.465 111.000 -60.155 113.515 ;
        RECT -63.015 101.145 -62.690 103.910 ;
        RECT -44.610 17.885 -44.250 204.515 ;
        RECT -26.845 130.910 -26.555 132.970 ;
        RECT -24.555 120.995 -24.230 123.760 ;
        RECT -17.975 121.120 -17.685 132.955 ;
        RECT -10.070 130.850 -9.760 133.365 ;
        RECT -12.620 120.995 -12.295 123.760 ;
        RECT 151.560 17.895 151.920 204.525 ;
        RECT 169.255 111.150 169.545 113.210 ;
        RECT 171.545 101.235 171.870 104.000 ;
        RECT 178.125 101.360 178.415 113.195 ;
        RECT 186.030 111.090 186.340 113.605 ;
        RECT 183.480 101.235 183.805 104.000 ;
        RECT 347.950 17.855 348.310 204.485 ;
        RECT 365.645 111.110 365.935 113.170 ;
        RECT 367.935 101.195 368.260 103.960 ;
        RECT 374.515 101.320 374.805 113.155 ;
        RECT 382.420 111.050 382.730 113.565 ;
        RECT 379.870 101.195 380.195 103.960 ;
        RECT 544.270 17.900 544.630 204.530 ;
        RECT 561.965 111.155 562.255 113.215 ;
        RECT 564.255 101.240 564.580 104.005 ;
        RECT 570.835 101.365 571.125 113.200 ;
        RECT 578.740 111.095 579.050 113.610 ;
        RECT 576.190 101.240 576.515 104.005 ;
        RECT 740.635 17.905 740.995 204.535 ;
        RECT 758.330 111.160 758.620 113.220 ;
        RECT 760.620 101.245 760.945 104.010 ;
        RECT 767.200 101.370 767.490 113.205 ;
        RECT 775.105 111.100 775.415 113.615 ;
        RECT 772.555 101.245 772.880 104.010 ;
        RECT 937.020 17.890 937.380 204.520 ;
        RECT 954.715 111.145 955.005 113.205 ;
        RECT 957.005 101.230 957.330 103.995 ;
        RECT 963.585 101.355 963.875 113.190 ;
        RECT 971.490 111.085 971.800 113.600 ;
        RECT 968.940 101.230 969.265 103.995 ;
        RECT 1133.345 17.895 1133.705 204.525 ;
        RECT 1151.040 111.150 1151.330 113.210 ;
        RECT 1153.330 101.235 1153.655 104.000 ;
        RECT 1159.910 101.360 1160.200 113.195 ;
        RECT 1167.815 111.090 1168.125 113.605 ;
        RECT 1165.265 101.235 1165.590 104.000 ;
    END
  END b6_p3
  PIN b7_q0
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT 1123.860 204.210 1125.480 204.535 ;
        RECT 1148.735 168.225 1149.115 168.605 ;
        RECT 1170.235 168.225 1170.615 168.605 ;
        RECT 1145.590 165.880 1164.260 165.890 ;
        RECT 1124.675 165.570 1172.245 165.880 ;
        RECT 1124.675 165.555 1145.885 165.570 ;
        RECT 1156.735 163.110 1157.115 163.115 ;
        RECT 1154.255 162.745 1157.120 163.110 ;
        RECT 1162.235 163.090 1162.615 163.115 ;
        RECT 1162.220 162.770 1164.365 163.090 ;
        RECT 1156.735 162.735 1157.115 162.745 ;
        RECT 1162.235 162.735 1162.615 162.770 ;
        RECT 1148.650 148.510 1149.030 148.890 ;
        RECT 1170.150 148.510 1170.530 148.890 ;
        RECT 1124.695 146.175 1145.715 146.185 ;
        RECT 1124.695 146.165 1164.175 146.175 ;
        RECT 1124.695 145.860 1172.160 146.165 ;
        RECT 1145.505 145.855 1172.160 145.860 ;
        RECT 1156.650 143.395 1157.030 143.400 ;
        RECT 1154.170 143.030 1157.035 143.395 ;
        RECT 1162.150 143.375 1162.530 143.400 ;
        RECT 1162.135 143.055 1164.280 143.375 ;
        RECT 1156.650 143.020 1157.030 143.030 ;
        RECT 1162.150 143.020 1162.530 143.055 ;
        RECT 1148.710 128.705 1149.090 129.085 ;
        RECT 1170.210 128.705 1170.590 129.085 ;
        RECT 1124.645 126.370 1145.925 126.375 ;
        RECT 1124.645 126.360 1164.235 126.370 ;
        RECT 1124.645 126.050 1172.220 126.360 ;
        RECT 1156.710 123.590 1157.090 123.595 ;
        RECT 1154.230 123.225 1157.095 123.590 ;
        RECT 1162.210 123.570 1162.590 123.595 ;
        RECT 1162.195 123.250 1164.340 123.570 ;
        RECT 1156.710 123.215 1157.090 123.225 ;
        RECT 1162.210 123.215 1162.590 123.250 ;
        RECT 1148.640 108.935 1149.020 109.315 ;
        RECT 1170.140 108.935 1170.520 109.315 ;
        RECT 1124.650 106.600 1145.695 106.615 ;
        RECT 1124.650 106.590 1164.165 106.600 ;
        RECT 1124.650 106.290 1172.150 106.590 ;
        RECT 1145.495 106.280 1172.150 106.290 ;
        RECT 1156.640 103.820 1157.020 103.825 ;
        RECT 1154.160 103.455 1157.025 103.820 ;
        RECT 1162.140 103.800 1162.520 103.825 ;
        RECT 1162.125 103.480 1164.270 103.800 ;
        RECT 1156.640 103.445 1157.020 103.455 ;
        RECT 1162.140 103.445 1162.520 103.480 ;
        RECT 1148.670 89.210 1149.050 89.590 ;
        RECT 1170.170 89.210 1170.550 89.590 ;
        RECT 1124.635 86.875 1145.715 86.880 ;
        RECT 1124.635 86.865 1164.195 86.875 ;
        RECT 1124.635 86.555 1172.180 86.865 ;
        RECT 1156.670 84.095 1157.050 84.100 ;
        RECT 1154.190 83.730 1157.055 84.095 ;
        RECT 1162.170 84.075 1162.550 84.100 ;
        RECT 1162.155 83.755 1164.300 84.075 ;
        RECT 1156.670 83.720 1157.050 83.730 ;
        RECT 1162.170 83.720 1162.550 83.755 ;
        RECT 1148.600 69.380 1148.980 69.760 ;
        RECT 1170.100 69.380 1170.480 69.760 ;
        RECT 1124.620 67.035 1164.125 67.045 ;
        RECT 1124.620 66.725 1172.110 67.035 ;
        RECT 1124.620 66.720 1145.640 66.725 ;
        RECT 1156.600 64.265 1156.980 64.270 ;
        RECT 1154.120 63.900 1156.985 64.265 ;
        RECT 1162.100 64.245 1162.480 64.270 ;
        RECT 1162.085 63.925 1164.230 64.245 ;
        RECT 1156.600 63.890 1156.980 63.900 ;
        RECT 1162.100 63.890 1162.480 63.925 ;
        RECT 1148.670 49.660 1149.050 50.040 ;
        RECT 1170.170 49.660 1170.550 50.040 ;
        RECT 1124.730 47.325 1145.780 47.335 ;
        RECT 1124.730 47.315 1164.195 47.325 ;
        RECT 1124.730 47.010 1172.180 47.315 ;
        RECT 1145.525 47.005 1172.180 47.010 ;
        RECT 1156.670 44.545 1157.050 44.550 ;
        RECT 1154.190 44.180 1157.055 44.545 ;
        RECT 1162.170 44.525 1162.550 44.550 ;
        RECT 1162.155 44.205 1164.300 44.525 ;
        RECT 1156.670 44.170 1157.050 44.180 ;
        RECT 1162.170 44.170 1162.550 44.205 ;
        RECT 1148.645 29.930 1149.025 30.310 ;
        RECT 1170.145 29.930 1170.525 30.310 ;
        RECT 1145.500 27.590 1164.170 27.595 ;
        RECT 1124.665 27.585 1164.170 27.590 ;
        RECT 1124.665 27.275 1172.155 27.585 ;
        RECT 1124.665 27.265 1145.645 27.275 ;
        RECT 1156.645 24.815 1157.025 24.820 ;
        RECT 1154.165 24.450 1157.030 24.815 ;
        RECT 1162.145 24.795 1162.525 24.820 ;
        RECT 1162.130 24.475 1164.275 24.795 ;
        RECT 1156.645 24.440 1157.025 24.450 ;
        RECT 1162.145 24.440 1162.525 24.475 ;
      LAYER Metal2 ;
        RECT 1124.885 17.840 1125.280 204.535 ;
        RECT 1148.685 165.570 1149.135 168.560 ;
        RECT 1154.410 162.560 1154.815 165.890 ;
        RECT 1163.845 162.615 1164.295 165.890 ;
        RECT 1170.200 165.570 1170.650 168.580 ;
        RECT 1148.600 145.855 1149.050 148.845 ;
        RECT 1154.325 142.845 1154.730 146.175 ;
        RECT 1163.760 142.900 1164.210 146.175 ;
        RECT 1170.115 145.855 1170.565 148.865 ;
        RECT 1148.660 126.050 1149.110 129.040 ;
        RECT 1154.385 123.040 1154.790 126.370 ;
        RECT 1163.820 123.095 1164.270 126.370 ;
        RECT 1170.175 126.050 1170.625 129.060 ;
        RECT 1148.590 106.280 1149.040 109.270 ;
        RECT 1154.315 103.270 1154.720 106.600 ;
        RECT 1163.750 103.325 1164.200 106.600 ;
        RECT 1170.105 106.280 1170.555 109.290 ;
        RECT 1148.620 86.555 1149.070 89.545 ;
        RECT 1154.345 83.545 1154.750 86.875 ;
        RECT 1163.780 83.600 1164.230 86.875 ;
        RECT 1170.135 86.555 1170.585 89.565 ;
        RECT 1148.550 66.725 1149.000 69.715 ;
        RECT 1154.275 63.715 1154.680 67.045 ;
        RECT 1163.710 63.770 1164.160 67.045 ;
        RECT 1170.065 66.725 1170.515 69.735 ;
        RECT 1148.620 47.005 1149.070 49.995 ;
        RECT 1154.345 43.995 1154.750 47.325 ;
        RECT 1163.780 44.050 1164.230 47.325 ;
        RECT 1170.135 47.005 1170.585 50.015 ;
        RECT 1148.595 27.275 1149.045 30.265 ;
        RECT 1154.320 24.265 1154.725 27.595 ;
        RECT 1163.755 24.320 1164.205 27.595 ;
        RECT 1170.110 27.275 1170.560 30.285 ;
    END
  END b7_q0
  PIN b7_q0_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT 1123.845 203.635 1126.405 203.940 ;
        RECT 1152.735 168.225 1153.115 168.605 ;
        RECT 1166.235 168.225 1166.615 168.605 ;
        RECT 1145.590 164.890 1172.245 164.900 ;
        RECT 1125.835 164.630 1172.245 164.890 ;
        RECT 1125.835 164.620 1145.830 164.630 ;
        RECT 1148.735 163.080 1149.115 163.115 ;
        RECT 1170.235 163.095 1170.615 163.115 ;
        RECT 1148.470 162.770 1151.480 163.080 ;
        RECT 1167.770 162.775 1170.680 163.095 ;
        RECT 1148.735 162.735 1149.115 162.770 ;
        RECT 1170.235 162.735 1170.615 162.775 ;
        RECT 1152.650 148.510 1153.030 148.890 ;
        RECT 1166.150 148.510 1166.530 148.890 ;
        RECT 1125.855 145.185 1145.660 145.195 ;
        RECT 1125.855 144.925 1172.160 145.185 ;
        RECT 1145.505 144.915 1172.160 144.925 ;
        RECT 1148.650 143.365 1149.030 143.400 ;
        RECT 1170.150 143.380 1170.530 143.400 ;
        RECT 1148.385 143.055 1151.395 143.365 ;
        RECT 1167.685 143.060 1170.595 143.380 ;
        RECT 1148.650 143.020 1149.030 143.055 ;
        RECT 1170.150 143.020 1170.530 143.060 ;
        RECT 1152.710 128.705 1153.090 129.085 ;
        RECT 1166.210 128.705 1166.590 129.085 ;
        RECT 1125.805 125.380 1145.890 125.385 ;
        RECT 1125.805 125.115 1172.220 125.380 ;
        RECT 1145.565 125.110 1172.220 125.115 ;
        RECT 1148.710 123.560 1149.090 123.595 ;
        RECT 1170.210 123.575 1170.590 123.595 ;
        RECT 1148.445 123.250 1151.455 123.560 ;
        RECT 1167.745 123.255 1170.655 123.575 ;
        RECT 1148.710 123.215 1149.090 123.250 ;
        RECT 1170.210 123.215 1170.590 123.255 ;
        RECT 1152.640 108.935 1153.020 109.315 ;
        RECT 1166.140 108.935 1166.520 109.315 ;
        RECT 1125.810 105.610 1145.715 105.625 ;
        RECT 1125.810 105.355 1172.150 105.610 ;
        RECT 1145.495 105.340 1172.150 105.355 ;
        RECT 1148.640 103.790 1149.020 103.825 ;
        RECT 1170.140 103.805 1170.520 103.825 ;
        RECT 1148.375 103.480 1151.385 103.790 ;
        RECT 1167.675 103.485 1170.585 103.805 ;
        RECT 1148.640 103.445 1149.020 103.480 ;
        RECT 1170.140 103.445 1170.520 103.485 ;
        RECT 1152.670 89.210 1153.050 89.590 ;
        RECT 1166.170 89.210 1166.550 89.590 ;
        RECT 1125.795 85.885 1145.770 85.890 ;
        RECT 1125.795 85.620 1172.180 85.885 ;
        RECT 1145.525 85.615 1172.180 85.620 ;
        RECT 1148.670 84.065 1149.050 84.100 ;
        RECT 1170.170 84.080 1170.550 84.100 ;
        RECT 1148.405 83.755 1151.415 84.065 ;
        RECT 1167.705 83.760 1170.615 84.080 ;
        RECT 1148.670 83.720 1149.050 83.755 ;
        RECT 1170.170 83.720 1170.550 83.760 ;
        RECT 1152.600 69.380 1152.980 69.760 ;
        RECT 1166.100 69.380 1166.480 69.760 ;
        RECT 1125.775 65.785 1172.110 66.055 ;
        RECT 1148.600 64.235 1148.980 64.270 ;
        RECT 1170.100 64.250 1170.480 64.270 ;
        RECT 1148.335 63.925 1151.345 64.235 ;
        RECT 1167.635 63.930 1170.545 64.250 ;
        RECT 1148.600 63.890 1148.980 63.925 ;
        RECT 1170.100 63.890 1170.480 63.930 ;
        RECT 1152.670 49.660 1153.050 50.040 ;
        RECT 1166.170 49.660 1166.550 50.040 ;
        RECT 1125.890 46.335 1145.780 46.345 ;
        RECT 1125.890 46.075 1172.180 46.335 ;
        RECT 1145.525 46.065 1172.180 46.075 ;
        RECT 1148.670 44.515 1149.050 44.550 ;
        RECT 1170.170 44.530 1170.550 44.550 ;
        RECT 1148.405 44.205 1151.415 44.515 ;
        RECT 1167.705 44.210 1170.615 44.530 ;
        RECT 1148.670 44.170 1149.050 44.205 ;
        RECT 1170.170 44.170 1170.550 44.210 ;
        RECT 1152.645 29.930 1153.025 30.310 ;
        RECT 1166.145 29.930 1166.525 30.310 ;
        RECT 1145.500 26.600 1172.155 26.605 ;
        RECT 1125.825 26.335 1172.155 26.600 ;
        RECT 1125.825 26.330 1145.725 26.335 ;
        RECT 1148.645 24.785 1149.025 24.820 ;
        RECT 1170.145 24.800 1170.525 24.820 ;
        RECT 1148.380 24.475 1151.390 24.785 ;
        RECT 1167.680 24.480 1170.590 24.800 ;
        RECT 1148.645 24.440 1149.025 24.475 ;
        RECT 1170.145 24.440 1170.525 24.480 ;
      LAYER Metal2 ;
        RECT 1125.990 17.925 1126.330 204.525 ;
        RECT 1151.085 162.585 1151.380 164.955 ;
        RECT 1152.695 164.630 1153.145 168.595 ;
        RECT 1166.225 164.630 1166.625 168.570 ;
        RECT 1167.875 162.620 1168.290 165.010 ;
        RECT 1151.000 142.870 1151.295 145.240 ;
        RECT 1152.610 144.915 1153.060 148.880 ;
        RECT 1166.140 144.915 1166.540 148.855 ;
        RECT 1167.790 142.905 1168.205 145.295 ;
        RECT 1151.060 123.065 1151.355 125.435 ;
        RECT 1152.670 125.110 1153.120 129.075 ;
        RECT 1166.200 125.110 1166.600 129.050 ;
        RECT 1167.850 123.100 1168.265 125.490 ;
        RECT 1150.990 103.295 1151.285 105.665 ;
        RECT 1152.600 105.340 1153.050 109.305 ;
        RECT 1166.130 105.340 1166.530 109.280 ;
        RECT 1167.780 103.330 1168.195 105.720 ;
        RECT 1151.020 83.570 1151.315 85.940 ;
        RECT 1152.630 85.615 1153.080 89.580 ;
        RECT 1166.160 85.615 1166.560 89.555 ;
        RECT 1167.810 83.605 1168.225 85.995 ;
        RECT 1150.950 63.740 1151.245 66.110 ;
        RECT 1152.560 65.785 1153.010 69.750 ;
        RECT 1166.090 65.785 1166.490 69.725 ;
        RECT 1167.740 63.775 1168.155 66.165 ;
        RECT 1151.020 44.020 1151.315 46.390 ;
        RECT 1152.630 46.065 1153.080 50.030 ;
        RECT 1166.160 46.065 1166.560 50.005 ;
        RECT 1167.810 44.055 1168.225 46.445 ;
        RECT 1150.995 24.290 1151.290 26.660 ;
        RECT 1152.605 26.335 1153.055 30.300 ;
        RECT 1166.135 26.335 1166.535 30.275 ;
        RECT 1167.785 24.325 1168.200 26.715 ;
    END
  END b7_q0_not
  PIN b1_q3
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.700 204.215 -102.185 204.530 ;
        RECT -79.545 168.135 -79.165 168.515 ;
        RECT -58.045 168.135 -57.665 168.515 ;
        RECT -103.050 165.790 -64.020 165.800 ;
        RECT -103.050 165.480 -56.035 165.790 ;
        RECT -103.050 165.475 -82.300 165.480 ;
        RECT -71.545 163.020 -71.165 163.025 ;
        RECT -74.025 162.655 -71.160 163.020 ;
        RECT -66.045 163.000 -65.665 163.025 ;
        RECT -66.060 162.680 -63.915 163.000 ;
        RECT -71.545 162.645 -71.165 162.655 ;
        RECT -66.045 162.645 -65.665 162.680 ;
        RECT -79.630 148.420 -79.250 148.800 ;
        RECT -58.130 148.420 -57.750 148.800 ;
        RECT -103.015 146.075 -64.105 146.085 ;
        RECT -103.015 145.765 -56.120 146.075 ;
        RECT -103.015 145.760 -82.265 145.765 ;
        RECT -71.630 143.305 -71.250 143.310 ;
        RECT -74.110 142.940 -71.245 143.305 ;
        RECT -66.130 143.285 -65.750 143.310 ;
        RECT -66.145 142.965 -64.000 143.285 ;
        RECT -71.630 142.930 -71.250 142.940 ;
        RECT -66.130 142.930 -65.750 142.965 ;
        RECT -79.570 128.615 -79.190 128.995 ;
        RECT -58.070 128.615 -57.690 128.995 ;
        RECT -82.715 126.275 -64.045 126.280 ;
        RECT -103.065 126.270 -64.045 126.275 ;
        RECT -103.065 125.960 -56.060 126.270 ;
        RECT -103.065 125.950 -82.315 125.960 ;
        RECT -71.570 123.500 -71.190 123.505 ;
        RECT -74.050 123.135 -71.185 123.500 ;
        RECT -66.070 123.480 -65.690 123.505 ;
        RECT -66.085 123.160 -63.940 123.480 ;
        RECT -71.570 123.125 -71.190 123.135 ;
        RECT -66.070 123.125 -65.690 123.160 ;
        RECT -79.640 108.845 -79.260 109.225 ;
        RECT -58.140 108.845 -57.760 109.225 ;
        RECT -103.060 106.510 -82.310 106.515 ;
        RECT -103.060 106.500 -64.115 106.510 ;
        RECT -103.060 106.190 -56.130 106.500 ;
        RECT -71.640 103.730 -71.260 103.735 ;
        RECT -74.120 103.365 -71.255 103.730 ;
        RECT -66.140 103.710 -65.760 103.735 ;
        RECT -66.155 103.390 -64.010 103.710 ;
        RECT -71.640 103.355 -71.260 103.365 ;
        RECT -66.140 103.355 -65.760 103.390 ;
        RECT -79.610 89.120 -79.230 89.500 ;
        RECT -58.110 89.120 -57.730 89.500 ;
        RECT -82.755 86.780 -64.085 86.785 ;
        RECT -103.075 86.775 -64.085 86.780 ;
        RECT -103.075 86.465 -56.100 86.775 ;
        RECT -103.075 86.455 -82.325 86.465 ;
        RECT -71.610 84.005 -71.230 84.010 ;
        RECT -74.090 83.640 -71.225 84.005 ;
        RECT -66.110 83.985 -65.730 84.010 ;
        RECT -66.125 83.665 -63.980 83.985 ;
        RECT -71.610 83.630 -71.230 83.640 ;
        RECT -66.110 83.630 -65.730 83.665 ;
        RECT -79.680 69.290 -79.300 69.670 ;
        RECT -58.180 69.290 -57.800 69.670 ;
        RECT -103.095 66.955 -82.345 66.970 ;
        RECT -103.095 66.945 -64.155 66.955 ;
        RECT -103.095 66.645 -56.170 66.945 ;
        RECT -82.825 66.635 -56.170 66.645 ;
        RECT -71.680 64.175 -71.300 64.180 ;
        RECT -74.160 63.810 -71.295 64.175 ;
        RECT -66.180 64.155 -65.800 64.180 ;
        RECT -66.195 63.835 -64.050 64.155 ;
        RECT -71.680 63.800 -71.300 63.810 ;
        RECT -66.180 63.800 -65.800 63.835 ;
        RECT -79.610 49.570 -79.230 49.950 ;
        RECT -58.110 49.570 -57.730 49.950 ;
        RECT -102.980 47.225 -64.085 47.235 ;
        RECT -102.980 46.915 -56.100 47.225 ;
        RECT -102.980 46.910 -82.230 46.915 ;
        RECT -71.610 44.455 -71.230 44.460 ;
        RECT -74.090 44.090 -71.225 44.455 ;
        RECT -66.110 44.435 -65.730 44.460 ;
        RECT -66.125 44.115 -63.980 44.435 ;
        RECT -71.610 44.080 -71.230 44.090 ;
        RECT -66.110 44.080 -65.730 44.115 ;
        RECT -79.605 29.760 -79.225 30.140 ;
        RECT -58.105 29.760 -57.725 30.140 ;
        RECT -82.750 27.420 -64.080 27.425 ;
        RECT -102.975 27.415 -64.080 27.420 ;
        RECT -102.975 27.105 -56.095 27.415 ;
        RECT -102.975 27.095 -82.225 27.105 ;
        RECT -71.605 24.645 -71.225 24.650 ;
        RECT -74.085 24.280 -71.220 24.645 ;
        RECT -66.105 24.625 -65.725 24.650 ;
        RECT -66.120 24.305 -63.975 24.625 ;
        RECT -71.605 24.270 -71.225 24.280 ;
        RECT -66.105 24.270 -65.725 24.305 ;
      LAYER Metal2 ;
        RECT -102.830 18.025 -102.435 204.530 ;
        RECT -79.595 165.480 -79.145 168.470 ;
        RECT -73.870 162.470 -73.465 165.800 ;
        RECT -64.435 162.525 -63.985 165.800 ;
        RECT -58.080 165.480 -57.630 168.490 ;
        RECT -79.680 145.765 -79.230 148.755 ;
        RECT -73.955 142.755 -73.550 146.085 ;
        RECT -64.520 142.810 -64.070 146.085 ;
        RECT -58.165 145.765 -57.715 148.775 ;
        RECT -79.620 125.960 -79.170 128.950 ;
        RECT -73.895 122.950 -73.490 126.280 ;
        RECT -64.460 123.005 -64.010 126.280 ;
        RECT -58.105 125.960 -57.655 128.970 ;
        RECT -79.690 106.190 -79.240 109.180 ;
        RECT -73.965 103.180 -73.560 106.510 ;
        RECT -64.530 103.235 -64.080 106.510 ;
        RECT -58.175 106.190 -57.725 109.200 ;
        RECT -79.660 86.465 -79.210 89.455 ;
        RECT -73.935 83.455 -73.530 86.785 ;
        RECT -64.500 83.510 -64.050 86.785 ;
        RECT -58.145 86.465 -57.695 89.475 ;
        RECT -79.730 66.635 -79.280 69.625 ;
        RECT -74.005 63.625 -73.600 66.955 ;
        RECT -64.570 63.680 -64.120 66.955 ;
        RECT -58.215 66.635 -57.765 69.645 ;
        RECT -79.660 46.915 -79.210 49.905 ;
        RECT -73.935 43.905 -73.530 47.235 ;
        RECT -64.500 43.960 -64.050 47.235 ;
        RECT -58.145 46.915 -57.695 49.925 ;
        RECT -79.655 27.105 -79.205 30.095 ;
        RECT -73.930 24.095 -73.525 27.425 ;
        RECT -64.495 24.150 -64.045 27.425 ;
        RECT -58.140 27.105 -57.690 30.115 ;
    END
  END b1_q3
  PIN p6_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 1112.085 168.835 1112.465 169.215 ;
        RECT 1109.010 168.340 1111.635 168.750 ;
        RECT 1111.195 165.900 1118.895 166.175 ;
        RECT 1111.210 162.475 1112.520 162.795 ;
        RECT 1109.020 161.920 1109.400 162.300 ;
      LAYER Metal2 ;
        RECT 1109.060 161.830 1109.360 168.770 ;
        RECT 1111.270 162.405 1111.550 168.765 ;
        RECT 1112.120 162.405 1112.420 169.225 ;
    END
  END p6_not
  PIN p6
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 1105.185 168.845 1105.565 169.225 ;
        RECT 1102.510 168.420 1104.250 168.710 ;
        RECT 1103.865 163.825 1119.885 164.160 ;
        RECT 1103.835 162.505 1105.615 162.795 ;
        RECT 1102.565 161.890 1102.945 162.270 ;
      LAYER Metal2 ;
        RECT 1102.595 161.830 1102.895 168.760 ;
        RECT 1103.905 162.430 1104.205 168.780 ;
        RECT 1105.220 162.460 1105.515 169.285 ;
    END
  END p6
  PIN p7_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 1308.425 168.835 1308.805 169.215 ;
        RECT 1305.350 168.340 1307.975 168.750 ;
        RECT 1307.535 165.900 1315.235 166.175 ;
        RECT 1307.550 162.475 1308.860 162.795 ;
        RECT 1305.360 161.920 1305.740 162.300 ;
      LAYER Metal2 ;
        RECT 1305.400 161.830 1305.700 168.770 ;
        RECT 1307.610 162.405 1307.890 168.765 ;
        RECT 1308.460 162.405 1308.760 169.225 ;
    END
  END p7_not
  PIN p7
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 1301.525 168.845 1301.905 169.225 ;
        RECT 1298.850 168.420 1300.590 168.710 ;
        RECT 1300.205 163.825 1316.225 164.160 ;
        RECT 1300.175 162.505 1301.955 162.795 ;
        RECT 1298.905 161.890 1299.285 162.270 ;
      LAYER Metal2 ;
        RECT 1298.935 161.830 1299.235 168.760 ;
        RECT 1300.245 162.430 1300.545 168.780 ;
        RECT 1301.560 162.460 1301.855 169.285 ;
    END
  END p7
  PIN p8_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 1308.225 149.110 1308.605 149.490 ;
        RECT 1305.150 148.615 1307.775 149.025 ;
        RECT 1307.335 146.175 1315.035 146.450 ;
        RECT 1307.350 142.750 1308.660 143.070 ;
        RECT 1305.160 142.195 1305.540 142.575 ;
      LAYER Metal2 ;
        RECT 1305.200 142.105 1305.500 149.045 ;
        RECT 1307.410 142.680 1307.690 149.040 ;
        RECT 1308.260 142.680 1308.560 149.500 ;
    END
  END p8_not
  PIN p8
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 1301.325 149.120 1301.705 149.500 ;
        RECT 1298.650 148.695 1300.390 148.985 ;
        RECT 1300.005 144.100 1316.025 144.435 ;
        RECT 1299.975 142.780 1301.755 143.070 ;
        RECT 1298.705 142.165 1299.085 142.545 ;
      LAYER Metal2 ;
        RECT 1298.735 142.105 1299.035 149.035 ;
        RECT 1300.045 142.705 1300.345 149.055 ;
        RECT 1301.360 142.735 1301.655 149.560 ;
    END
  END p8
  PIN p9_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 1308.380 129.465 1308.760 129.845 ;
        RECT 1305.305 128.970 1307.930 129.380 ;
        RECT 1307.490 126.530 1315.190 126.805 ;
        RECT 1307.505 123.105 1308.815 123.425 ;
        RECT 1305.315 122.550 1305.695 122.930 ;
      LAYER Metal2 ;
        RECT 1305.355 122.460 1305.655 129.400 ;
        RECT 1307.565 123.035 1307.845 129.395 ;
        RECT 1308.415 123.035 1308.715 129.855 ;
    END
  END p9_not
  PIN p9
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 1301.480 129.475 1301.860 129.855 ;
        RECT 1298.805 129.050 1300.545 129.340 ;
        RECT 1300.160 124.455 1316.180 124.790 ;
        RECT 1300.130 123.135 1301.910 123.425 ;
        RECT 1298.860 122.520 1299.240 122.900 ;
      LAYER Metal2 ;
        RECT 1298.890 122.460 1299.190 129.390 ;
        RECT 1300.200 123.060 1300.500 129.410 ;
        RECT 1301.515 123.090 1301.810 129.915 ;
    END
  END p9
  PIN p10_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 1308.380 109.670 1308.760 110.050 ;
        RECT 1305.305 109.175 1307.930 109.585 ;
        RECT 1307.490 106.735 1315.190 107.010 ;
        RECT 1307.505 103.310 1308.815 103.630 ;
        RECT 1305.315 102.755 1305.695 103.135 ;
      LAYER Metal2 ;
        RECT 1305.355 102.665 1305.655 109.605 ;
        RECT 1307.565 103.240 1307.845 109.600 ;
        RECT 1308.415 103.240 1308.715 110.060 ;
    END
  END p10_not
  PIN p10
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 1301.480 109.680 1301.860 110.060 ;
        RECT 1298.805 109.255 1300.545 109.545 ;
        RECT 1300.160 104.660 1316.180 104.995 ;
        RECT 1300.130 103.340 1301.910 103.630 ;
        RECT 1298.860 102.725 1299.240 103.105 ;
      LAYER Metal2 ;
        RECT 1298.890 102.665 1299.190 109.595 ;
        RECT 1300.200 103.265 1300.500 109.615 ;
        RECT 1301.515 103.295 1301.810 110.120 ;
    END
  END p10
  PIN b7_c0_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1147.100 171.225 1148.555 171.605 ;
        RECT 1147.260 168.925 1148.555 169.305 ;
        RECT 1160.745 168.925 1162.055 169.305 ;
        RECT 1145.590 167.600 1161.600 167.975 ;
        RECT 1147.270 163.425 1148.575 163.805 ;
        RECT 1160.610 163.425 1162.075 163.805 ;
        RECT 1147.085 161.425 1148.575 161.805 ;
      LAYER Metal2 ;
        RECT 1147.390 160.715 1147.745 171.800 ;
        RECT 1160.900 163.145 1161.230 169.340 ;
    END
  END b7_c0_not
  PIN b7_c1_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1147.015 151.510 1148.470 151.890 ;
        RECT 1147.175 149.210 1148.470 149.590 ;
        RECT 1160.660 149.210 1161.970 149.590 ;
        RECT 1145.505 147.885 1161.515 148.260 ;
        RECT 1147.185 143.710 1148.490 144.090 ;
        RECT 1160.525 143.710 1161.990 144.090 ;
        RECT 1147.000 141.710 1148.490 142.090 ;
      LAYER Metal2 ;
        RECT 1147.305 141.000 1147.660 152.085 ;
        RECT 1160.815 143.430 1161.145 149.625 ;
    END
  END b7_c1_not
  PIN b7_c0
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1170.795 171.325 1172.075 171.705 ;
        RECT 1157.295 168.925 1158.480 169.305 ;
        RECT 1170.795 168.925 1171.810 169.305 ;
        RECT 1145.590 166.245 1171.820 166.635 ;
        RECT 1157.275 163.425 1158.635 163.805 ;
        RECT 1170.775 163.425 1171.955 163.805 ;
        RECT 1170.775 161.425 1171.850 161.805 ;
      LAYER Metal2 ;
        RECT 1157.915 169.290 1158.225 169.320 ;
        RECT 1157.915 163.190 1158.230 169.290 ;
        RECT 1171.415 161.195 1171.745 171.890 ;
    END
  END b7_c0
  PIN b7_c1
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1170.710 151.610 1171.990 151.990 ;
        RECT 1157.210 149.210 1158.395 149.590 ;
        RECT 1170.710 149.210 1171.725 149.590 ;
        RECT 1145.505 146.530 1171.735 146.920 ;
        RECT 1157.190 143.710 1158.550 144.090 ;
        RECT 1170.690 143.710 1171.870 144.090 ;
        RECT 1170.690 141.710 1171.765 142.090 ;
      LAYER Metal2 ;
        RECT 1157.830 149.575 1158.140 149.605 ;
        RECT 1157.830 143.475 1158.145 149.575 ;
        RECT 1171.330 141.480 1171.660 152.175 ;
    END
  END b7_c1
  PIN b7_c2_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1147.075 131.705 1148.530 132.085 ;
        RECT 1147.235 129.405 1148.530 129.785 ;
        RECT 1160.720 129.405 1162.030 129.785 ;
        RECT 1145.565 128.080 1161.575 128.455 ;
        RECT 1147.245 123.905 1148.550 124.285 ;
        RECT 1160.585 123.905 1162.050 124.285 ;
        RECT 1147.060 121.905 1148.550 122.285 ;
      LAYER Metal2 ;
        RECT 1147.365 121.195 1147.720 132.280 ;
        RECT 1160.875 123.625 1161.205 129.820 ;
    END
  END b7_c2_not
  PIN b7_c2
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1170.770 131.805 1172.050 132.185 ;
        RECT 1157.270 129.405 1158.455 129.785 ;
        RECT 1170.770 129.405 1171.785 129.785 ;
        RECT 1145.565 126.725 1171.795 127.115 ;
        RECT 1157.250 123.905 1158.610 124.285 ;
        RECT 1170.750 123.905 1171.930 124.285 ;
        RECT 1170.750 121.905 1171.825 122.285 ;
      LAYER Metal2 ;
        RECT 1157.890 129.770 1158.200 129.800 ;
        RECT 1157.890 123.670 1158.205 129.770 ;
        RECT 1171.390 121.675 1171.720 132.370 ;
    END
  END b7_c2
  PIN b7_c3_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1147.005 111.935 1148.460 112.315 ;
        RECT 1147.165 109.635 1148.460 110.015 ;
        RECT 1160.650 109.635 1161.960 110.015 ;
        RECT 1145.495 108.310 1161.505 108.685 ;
        RECT 1147.175 104.135 1148.480 104.515 ;
        RECT 1160.515 104.135 1161.980 104.515 ;
        RECT 1146.990 102.135 1148.480 102.515 ;
      LAYER Metal2 ;
        RECT 1147.295 101.425 1147.650 112.510 ;
        RECT 1160.805 103.855 1161.135 110.050 ;
    END
  END b7_c3_not
  PIN b7_c3
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1170.700 112.035 1171.980 112.415 ;
        RECT 1157.200 109.635 1158.385 110.015 ;
        RECT 1170.700 109.635 1171.715 110.015 ;
        RECT 1145.495 106.955 1171.725 107.345 ;
        RECT 1157.180 104.135 1158.540 104.515 ;
        RECT 1170.680 104.135 1171.860 104.515 ;
        RECT 1170.680 102.135 1171.755 102.515 ;
      LAYER Metal2 ;
        RECT 1157.820 110.000 1158.130 110.030 ;
        RECT 1157.820 103.900 1158.135 110.000 ;
        RECT 1171.320 101.905 1171.650 112.600 ;
    END
  END b7_c3
  PIN b5_c0
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 778.085 171.335 779.365 171.715 ;
        RECT 764.585 168.935 765.770 169.315 ;
        RECT 778.085 168.935 779.100 169.315 ;
        RECT 752.880 166.255 779.110 166.645 ;
        RECT 764.565 163.435 765.925 163.815 ;
        RECT 778.065 163.435 779.245 163.815 ;
        RECT 778.065 161.435 779.140 161.815 ;
      LAYER Metal2 ;
        RECT 765.205 169.300 765.515 169.330 ;
        RECT 765.205 163.200 765.520 169.300 ;
        RECT 778.705 161.205 779.035 171.900 ;
    END
  END b5_c0
  PIN b5_c0_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 754.390 171.235 755.845 171.615 ;
        RECT 754.550 168.935 755.845 169.315 ;
        RECT 768.035 168.935 769.345 169.315 ;
        RECT 752.880 167.610 768.890 167.985 ;
        RECT 754.560 163.435 755.865 163.815 ;
        RECT 767.900 163.435 769.365 163.815 ;
        RECT 754.375 161.435 755.865 161.815 ;
      LAYER Metal2 ;
        RECT 754.680 160.725 755.035 171.810 ;
        RECT 768.190 163.155 768.520 169.350 ;
    END
  END b5_c0_not
  PIN b5
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT 731.150 204.220 732.770 204.545 ;
        RECT 756.025 168.235 756.405 168.615 ;
        RECT 777.525 168.235 777.905 168.615 ;
        RECT 752.880 165.890 771.550 165.900 ;
        RECT 731.965 165.580 779.535 165.890 ;
        RECT 731.965 165.565 753.175 165.580 ;
        RECT 764.025 163.120 764.405 163.125 ;
        RECT 761.545 162.755 764.410 163.120 ;
        RECT 769.525 163.100 769.905 163.125 ;
        RECT 769.510 162.780 771.655 163.100 ;
        RECT 764.025 162.745 764.405 162.755 ;
        RECT 769.525 162.745 769.905 162.780 ;
        RECT 755.940 148.520 756.320 148.900 ;
        RECT 777.440 148.520 777.820 148.900 ;
        RECT 731.985 146.185 753.005 146.195 ;
        RECT 731.985 146.175 771.465 146.185 ;
        RECT 731.985 145.870 779.450 146.175 ;
        RECT 752.795 145.865 779.450 145.870 ;
        RECT 763.940 143.405 764.320 143.410 ;
        RECT 761.460 143.040 764.325 143.405 ;
        RECT 769.440 143.385 769.820 143.410 ;
        RECT 769.425 143.065 771.570 143.385 ;
        RECT 763.940 143.030 764.320 143.040 ;
        RECT 769.440 143.030 769.820 143.065 ;
        RECT 756.000 128.715 756.380 129.095 ;
        RECT 777.500 128.715 777.880 129.095 ;
        RECT 731.935 126.380 753.215 126.385 ;
        RECT 731.935 126.370 771.525 126.380 ;
        RECT 731.935 126.060 779.510 126.370 ;
        RECT 764.000 123.600 764.380 123.605 ;
        RECT 761.520 123.235 764.385 123.600 ;
        RECT 769.500 123.580 769.880 123.605 ;
        RECT 769.485 123.260 771.630 123.580 ;
        RECT 764.000 123.225 764.380 123.235 ;
        RECT 769.500 123.225 769.880 123.260 ;
        RECT 755.930 108.945 756.310 109.325 ;
        RECT 777.430 108.945 777.810 109.325 ;
        RECT 731.940 106.610 752.985 106.625 ;
        RECT 731.940 106.600 771.455 106.610 ;
        RECT 731.940 106.300 779.440 106.600 ;
        RECT 752.785 106.290 779.440 106.300 ;
        RECT 763.930 103.830 764.310 103.835 ;
        RECT 761.450 103.465 764.315 103.830 ;
        RECT 769.430 103.810 769.810 103.835 ;
        RECT 769.415 103.490 771.560 103.810 ;
        RECT 763.930 103.455 764.310 103.465 ;
        RECT 769.430 103.455 769.810 103.490 ;
        RECT 755.960 89.220 756.340 89.600 ;
        RECT 777.460 89.220 777.840 89.600 ;
        RECT 731.925 86.885 753.005 86.890 ;
        RECT 731.925 86.875 771.485 86.885 ;
        RECT 731.925 86.565 779.470 86.875 ;
        RECT 763.960 84.105 764.340 84.110 ;
        RECT 761.480 83.740 764.345 84.105 ;
        RECT 769.460 84.085 769.840 84.110 ;
        RECT 769.445 83.765 771.590 84.085 ;
        RECT 763.960 83.730 764.340 83.740 ;
        RECT 769.460 83.730 769.840 83.765 ;
        RECT 755.890 69.390 756.270 69.770 ;
        RECT 777.390 69.390 777.770 69.770 ;
        RECT 731.910 67.045 771.415 67.055 ;
        RECT 731.910 66.735 779.400 67.045 ;
        RECT 731.910 66.730 752.930 66.735 ;
        RECT 763.890 64.275 764.270 64.280 ;
        RECT 761.410 63.910 764.275 64.275 ;
        RECT 769.390 64.255 769.770 64.280 ;
        RECT 769.375 63.935 771.520 64.255 ;
        RECT 763.890 63.900 764.270 63.910 ;
        RECT 769.390 63.900 769.770 63.935 ;
        RECT 755.960 49.670 756.340 50.050 ;
        RECT 777.460 49.670 777.840 50.050 ;
        RECT 732.020 47.335 753.070 47.345 ;
        RECT 732.020 47.325 771.485 47.335 ;
        RECT 732.020 47.020 779.470 47.325 ;
        RECT 752.815 47.015 779.470 47.020 ;
        RECT 763.960 44.555 764.340 44.560 ;
        RECT 761.480 44.190 764.345 44.555 ;
        RECT 769.460 44.535 769.840 44.560 ;
        RECT 769.445 44.215 771.590 44.535 ;
        RECT 763.960 44.180 764.340 44.190 ;
        RECT 769.460 44.180 769.840 44.215 ;
        RECT 755.935 29.940 756.315 30.320 ;
        RECT 777.435 29.940 777.815 30.320 ;
        RECT 752.790 27.600 771.460 27.605 ;
        RECT 731.955 27.595 771.460 27.600 ;
        RECT 731.955 27.285 779.445 27.595 ;
        RECT 731.955 27.275 752.935 27.285 ;
        RECT 763.935 24.825 764.315 24.830 ;
        RECT 761.455 24.460 764.320 24.825 ;
        RECT 769.435 24.805 769.815 24.830 ;
        RECT 769.420 24.485 771.565 24.805 ;
        RECT 763.935 24.450 764.315 24.460 ;
        RECT 769.435 24.450 769.815 24.485 ;
      LAYER Metal2 ;
        RECT 732.175 17.850 732.570 204.545 ;
        RECT 755.975 165.580 756.425 168.570 ;
        RECT 761.700 162.570 762.105 165.900 ;
        RECT 771.135 162.625 771.585 165.900 ;
        RECT 777.490 165.580 777.940 168.590 ;
        RECT 755.890 145.865 756.340 148.855 ;
        RECT 761.615 142.855 762.020 146.185 ;
        RECT 771.050 142.910 771.500 146.185 ;
        RECT 777.405 145.865 777.855 148.875 ;
        RECT 755.950 126.060 756.400 129.050 ;
        RECT 761.675 123.050 762.080 126.380 ;
        RECT 771.110 123.105 771.560 126.380 ;
        RECT 777.465 126.060 777.915 129.070 ;
        RECT 755.880 106.290 756.330 109.280 ;
        RECT 761.605 103.280 762.010 106.610 ;
        RECT 771.040 103.335 771.490 106.610 ;
        RECT 777.395 106.290 777.845 109.300 ;
        RECT 755.910 86.565 756.360 89.555 ;
        RECT 761.635 83.555 762.040 86.885 ;
        RECT 771.070 83.610 771.520 86.885 ;
        RECT 777.425 86.565 777.875 89.575 ;
        RECT 755.840 66.735 756.290 69.725 ;
        RECT 761.565 63.725 761.970 67.055 ;
        RECT 771.000 63.780 771.450 67.055 ;
        RECT 777.355 66.735 777.805 69.745 ;
        RECT 755.910 47.015 756.360 50.005 ;
        RECT 761.635 44.005 762.040 47.335 ;
        RECT 771.070 44.060 771.520 47.335 ;
        RECT 777.425 47.015 777.875 50.025 ;
        RECT 755.885 27.285 756.335 30.275 ;
        RECT 761.610 24.275 762.015 27.605 ;
        RECT 771.045 24.330 771.495 27.605 ;
        RECT 777.400 27.285 777.850 30.295 ;
    END
  END b5
  PIN b5_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT 731.135 203.645 733.695 203.950 ;
        RECT 760.025 168.235 760.405 168.615 ;
        RECT 773.525 168.235 773.905 168.615 ;
        RECT 752.880 164.900 779.535 164.910 ;
        RECT 733.125 164.640 779.535 164.900 ;
        RECT 733.125 164.630 753.120 164.640 ;
        RECT 756.025 163.090 756.405 163.125 ;
        RECT 777.525 163.105 777.905 163.125 ;
        RECT 755.760 162.780 758.770 163.090 ;
        RECT 775.060 162.785 777.970 163.105 ;
        RECT 756.025 162.745 756.405 162.780 ;
        RECT 777.525 162.745 777.905 162.785 ;
        RECT 759.940 148.520 760.320 148.900 ;
        RECT 773.440 148.520 773.820 148.900 ;
        RECT 733.145 145.195 752.950 145.205 ;
        RECT 733.145 144.935 779.450 145.195 ;
        RECT 752.795 144.925 779.450 144.935 ;
        RECT 755.940 143.375 756.320 143.410 ;
        RECT 777.440 143.390 777.820 143.410 ;
        RECT 755.675 143.065 758.685 143.375 ;
        RECT 774.975 143.070 777.885 143.390 ;
        RECT 755.940 143.030 756.320 143.065 ;
        RECT 777.440 143.030 777.820 143.070 ;
        RECT 760.000 128.715 760.380 129.095 ;
        RECT 773.500 128.715 773.880 129.095 ;
        RECT 733.095 125.390 753.180 125.395 ;
        RECT 733.095 125.125 779.510 125.390 ;
        RECT 752.855 125.120 779.510 125.125 ;
        RECT 756.000 123.570 756.380 123.605 ;
        RECT 777.500 123.585 777.880 123.605 ;
        RECT 755.735 123.260 758.745 123.570 ;
        RECT 775.035 123.265 777.945 123.585 ;
        RECT 756.000 123.225 756.380 123.260 ;
        RECT 777.500 123.225 777.880 123.265 ;
        RECT 759.930 108.945 760.310 109.325 ;
        RECT 773.430 108.945 773.810 109.325 ;
        RECT 733.100 105.620 753.005 105.635 ;
        RECT 733.100 105.365 779.440 105.620 ;
        RECT 752.785 105.350 779.440 105.365 ;
        RECT 755.930 103.800 756.310 103.835 ;
        RECT 777.430 103.815 777.810 103.835 ;
        RECT 755.665 103.490 758.675 103.800 ;
        RECT 774.965 103.495 777.875 103.815 ;
        RECT 755.930 103.455 756.310 103.490 ;
        RECT 777.430 103.455 777.810 103.495 ;
        RECT 759.960 89.220 760.340 89.600 ;
        RECT 773.460 89.220 773.840 89.600 ;
        RECT 733.085 85.895 753.060 85.900 ;
        RECT 733.085 85.630 779.470 85.895 ;
        RECT 752.815 85.625 779.470 85.630 ;
        RECT 755.960 84.075 756.340 84.110 ;
        RECT 777.460 84.090 777.840 84.110 ;
        RECT 755.695 83.765 758.705 84.075 ;
        RECT 774.995 83.770 777.905 84.090 ;
        RECT 755.960 83.730 756.340 83.765 ;
        RECT 777.460 83.730 777.840 83.770 ;
        RECT 759.890 69.390 760.270 69.770 ;
        RECT 773.390 69.390 773.770 69.770 ;
        RECT 733.065 65.795 779.400 66.065 ;
        RECT 755.890 64.245 756.270 64.280 ;
        RECT 777.390 64.260 777.770 64.280 ;
        RECT 755.625 63.935 758.635 64.245 ;
        RECT 774.925 63.940 777.835 64.260 ;
        RECT 755.890 63.900 756.270 63.935 ;
        RECT 777.390 63.900 777.770 63.940 ;
        RECT 759.960 49.670 760.340 50.050 ;
        RECT 773.460 49.670 773.840 50.050 ;
        RECT 733.180 46.345 753.070 46.355 ;
        RECT 733.180 46.085 779.470 46.345 ;
        RECT 752.815 46.075 779.470 46.085 ;
        RECT 755.960 44.525 756.340 44.560 ;
        RECT 777.460 44.540 777.840 44.560 ;
        RECT 755.695 44.215 758.705 44.525 ;
        RECT 774.995 44.220 777.905 44.540 ;
        RECT 755.960 44.180 756.340 44.215 ;
        RECT 777.460 44.180 777.840 44.220 ;
        RECT 759.935 29.940 760.315 30.320 ;
        RECT 773.435 29.940 773.815 30.320 ;
        RECT 752.790 26.610 779.445 26.615 ;
        RECT 733.115 26.345 779.445 26.610 ;
        RECT 733.115 26.340 753.015 26.345 ;
        RECT 755.935 24.795 756.315 24.830 ;
        RECT 777.435 24.810 777.815 24.830 ;
        RECT 755.670 24.485 758.680 24.795 ;
        RECT 774.970 24.490 777.880 24.810 ;
        RECT 755.935 24.450 756.315 24.485 ;
        RECT 777.435 24.450 777.815 24.490 ;
      LAYER Metal2 ;
        RECT 733.280 17.935 733.620 204.535 ;
        RECT 758.375 162.595 758.670 164.965 ;
        RECT 759.985 164.640 760.435 168.605 ;
        RECT 773.515 164.640 773.915 168.580 ;
        RECT 775.165 162.630 775.580 165.020 ;
        RECT 758.290 142.880 758.585 145.250 ;
        RECT 759.900 144.925 760.350 148.890 ;
        RECT 773.430 144.925 773.830 148.865 ;
        RECT 775.080 142.915 775.495 145.305 ;
        RECT 758.350 123.075 758.645 125.445 ;
        RECT 759.960 125.120 760.410 129.085 ;
        RECT 773.490 125.120 773.890 129.060 ;
        RECT 775.140 123.110 775.555 125.500 ;
        RECT 758.280 103.305 758.575 105.675 ;
        RECT 759.890 105.350 760.340 109.315 ;
        RECT 773.420 105.350 773.820 109.290 ;
        RECT 775.070 103.340 775.485 105.730 ;
        RECT 758.310 83.580 758.605 85.950 ;
        RECT 759.920 85.625 760.370 89.590 ;
        RECT 773.450 85.625 773.850 89.565 ;
        RECT 775.100 83.615 775.515 86.005 ;
        RECT 758.240 63.750 758.535 66.120 ;
        RECT 759.850 65.795 760.300 69.760 ;
        RECT 773.380 65.795 773.780 69.735 ;
        RECT 775.030 63.785 775.445 66.175 ;
        RECT 758.310 44.030 758.605 46.400 ;
        RECT 759.920 46.075 760.370 50.040 ;
        RECT 773.450 46.075 773.850 50.015 ;
        RECT 775.100 44.065 775.515 46.455 ;
        RECT 758.285 24.300 758.580 26.670 ;
        RECT 759.895 26.345 760.345 30.310 ;
        RECT 773.425 26.345 773.825 30.285 ;
        RECT 775.075 24.335 775.490 26.725 ;
    END
  END b5_not
  PIN p4_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 719.405 168.835 719.785 169.215 ;
        RECT 716.330 168.340 718.955 168.750 ;
        RECT 718.515 165.900 726.215 166.175 ;
        RECT 718.530 162.475 719.840 162.795 ;
        RECT 716.340 161.920 716.720 162.300 ;
      LAYER Metal2 ;
        RECT 716.380 161.830 716.680 168.770 ;
        RECT 718.590 162.405 718.870 168.765 ;
        RECT 719.440 162.405 719.740 169.225 ;
    END
  END p4_not
  PIN p4
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 712.505 168.845 712.885 169.225 ;
        RECT 709.830 168.420 711.570 168.710 ;
        RECT 711.185 163.825 727.205 164.160 ;
        RECT 711.155 162.505 712.935 162.795 ;
        RECT 709.885 161.890 710.265 162.270 ;
      LAYER Metal2 ;
        RECT 709.915 161.830 710.215 168.760 ;
        RECT 711.225 162.430 711.525 168.780 ;
        RECT 712.540 162.460 712.835 169.285 ;
    END
  END p4
  PIN p5_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 915.745 168.835 916.125 169.215 ;
        RECT 912.670 168.340 915.295 168.750 ;
        RECT 914.855 165.900 922.555 166.175 ;
        RECT 914.870 162.475 916.180 162.795 ;
        RECT 912.680 161.920 913.060 162.300 ;
      LAYER Metal2 ;
        RECT 912.720 161.830 913.020 168.770 ;
        RECT 914.930 162.405 915.210 168.765 ;
        RECT 915.780 162.405 916.080 169.225 ;
    END
  END p5_not
  PIN p5
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 908.845 168.845 909.225 169.225 ;
        RECT 906.170 168.420 907.910 168.710 ;
        RECT 907.525 163.825 923.545 164.160 ;
        RECT 907.495 162.505 909.275 162.795 ;
        RECT 906.225 161.890 906.605 162.270 ;
      LAYER Metal2 ;
        RECT 906.255 161.830 906.555 168.760 ;
        RECT 907.565 162.430 907.865 168.780 ;
        RECT 908.880 162.460 909.175 169.285 ;
    END
  END p5
  PIN b5_c2_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 754.365 131.715 755.820 132.095 ;
        RECT 754.525 129.415 755.820 129.795 ;
        RECT 768.010 129.415 769.320 129.795 ;
        RECT 752.855 128.090 768.865 128.465 ;
        RECT 754.535 123.915 755.840 124.295 ;
        RECT 767.875 123.915 769.340 124.295 ;
        RECT 754.350 121.915 755.840 122.295 ;
      LAYER Metal2 ;
        RECT 754.655 121.205 755.010 132.290 ;
        RECT 768.165 123.635 768.495 129.830 ;
    END
  END b5_c2_not
  PIN b6_c0_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 950.775 171.220 952.230 171.600 ;
        RECT 950.935 168.920 952.230 169.300 ;
        RECT 964.420 168.920 965.730 169.300 ;
        RECT 949.265 167.595 965.275 167.970 ;
        RECT 950.945 163.420 952.250 163.800 ;
        RECT 964.285 163.420 965.750 163.800 ;
        RECT 950.760 161.420 952.250 161.800 ;
      LAYER Metal2 ;
        RECT 951.065 160.710 951.420 171.795 ;
        RECT 964.575 163.140 964.905 169.335 ;
    END
  END b6_c0_not
  PIN b6_c1_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 950.690 151.505 952.145 151.885 ;
        RECT 950.850 149.205 952.145 149.585 ;
        RECT 964.335 149.205 965.645 149.585 ;
        RECT 949.180 147.880 965.190 148.255 ;
        RECT 950.860 143.705 952.165 144.085 ;
        RECT 964.200 143.705 965.665 144.085 ;
        RECT 950.675 141.705 952.165 142.085 ;
      LAYER Metal2 ;
        RECT 950.980 140.995 951.335 152.080 ;
        RECT 964.490 143.425 964.820 149.620 ;
    END
  END b6_c1_not
  PIN b6_c0
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 974.470 171.320 975.750 171.700 ;
        RECT 960.970 168.920 962.155 169.300 ;
        RECT 974.470 168.920 975.485 169.300 ;
        RECT 949.265 166.240 975.495 166.630 ;
        RECT 960.950 163.420 962.310 163.800 ;
        RECT 974.450 163.420 975.630 163.800 ;
        RECT 974.450 161.420 975.525 161.800 ;
      LAYER Metal2 ;
        RECT 961.590 169.285 961.900 169.315 ;
        RECT 961.590 163.185 961.905 169.285 ;
        RECT 975.090 161.190 975.420 171.885 ;
    END
  END b6_c0
  PIN b6_c1
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 974.385 151.605 975.665 151.985 ;
        RECT 960.885 149.205 962.070 149.585 ;
        RECT 974.385 149.205 975.400 149.585 ;
        RECT 949.180 146.525 975.410 146.915 ;
        RECT 960.865 143.705 962.225 144.085 ;
        RECT 974.365 143.705 975.545 144.085 ;
        RECT 974.365 141.705 975.440 142.085 ;
      LAYER Metal2 ;
        RECT 961.505 149.570 961.815 149.600 ;
        RECT 961.505 143.470 961.820 149.570 ;
        RECT 975.005 141.475 975.335 152.170 ;
    END
  END b6_c1
  PIN b6_c2_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 950.750 131.700 952.205 132.080 ;
        RECT 950.910 129.400 952.205 129.780 ;
        RECT 964.395 129.400 965.705 129.780 ;
        RECT 949.240 128.075 965.250 128.450 ;
        RECT 950.920 123.900 952.225 124.280 ;
        RECT 964.260 123.900 965.725 124.280 ;
        RECT 950.735 121.900 952.225 122.280 ;
      LAYER Metal2 ;
        RECT 951.040 121.190 951.395 132.275 ;
        RECT 964.550 123.620 964.880 129.815 ;
    END
  END b6_c2_not
  PIN b6_c2
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 974.445 131.800 975.725 132.180 ;
        RECT 960.945 129.400 962.130 129.780 ;
        RECT 974.445 129.400 975.460 129.780 ;
        RECT 949.240 126.720 975.470 127.110 ;
        RECT 960.925 123.900 962.285 124.280 ;
        RECT 974.425 123.900 975.605 124.280 ;
        RECT 974.425 121.900 975.500 122.280 ;
      LAYER Metal2 ;
        RECT 961.565 129.765 961.875 129.795 ;
        RECT 961.565 123.665 961.880 129.765 ;
        RECT 975.065 121.670 975.395 132.365 ;
    END
  END b6_c2
  PIN b6_c3_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 950.680 111.930 952.135 112.310 ;
        RECT 950.840 109.630 952.135 110.010 ;
        RECT 964.325 109.630 965.635 110.010 ;
        RECT 949.170 108.305 965.180 108.680 ;
        RECT 950.850 104.130 952.155 104.510 ;
        RECT 964.190 104.130 965.655 104.510 ;
        RECT 950.665 102.130 952.155 102.510 ;
      LAYER Metal2 ;
        RECT 950.970 101.420 951.325 112.505 ;
        RECT 964.480 103.850 964.810 110.045 ;
    END
  END b6_c3_not
  PIN b6_c3
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 974.375 112.030 975.655 112.410 ;
        RECT 960.875 109.630 962.060 110.010 ;
        RECT 974.375 109.630 975.390 110.010 ;
        RECT 949.170 106.950 975.400 107.340 ;
        RECT 960.855 104.130 962.215 104.510 ;
        RECT 974.355 104.130 975.535 104.510 ;
        RECT 974.355 102.130 975.430 102.510 ;
      LAYER Metal2 ;
        RECT 961.495 109.995 961.805 110.025 ;
        RECT 961.495 103.895 961.810 109.995 ;
        RECT 974.995 101.900 975.325 112.595 ;
    END
  END b6_c3
  PIN b5_c3
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 777.990 112.045 779.270 112.425 ;
        RECT 764.490 109.645 765.675 110.025 ;
        RECT 777.990 109.645 779.005 110.025 ;
        RECT 752.785 106.965 779.015 107.355 ;
        RECT 764.470 104.145 765.830 104.525 ;
        RECT 777.970 104.145 779.150 104.525 ;
        RECT 777.970 102.145 779.045 102.525 ;
      LAYER Metal2 ;
        RECT 765.110 110.010 765.420 110.040 ;
        RECT 765.110 103.910 765.425 110.010 ;
        RECT 778.610 101.915 778.940 112.610 ;
    END
  END b5_c3
  PIN b5_c3_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 754.295 111.945 755.750 112.325 ;
        RECT 754.455 109.645 755.750 110.025 ;
        RECT 767.940 109.645 769.250 110.025 ;
        RECT 752.785 108.320 768.795 108.695 ;
        RECT 754.465 104.145 755.770 104.525 ;
        RECT 767.805 104.145 769.270 104.525 ;
        RECT 754.280 102.145 755.770 102.525 ;
      LAYER Metal2 ;
        RECT 754.585 101.435 754.940 112.520 ;
        RECT 768.095 103.865 768.425 110.060 ;
    END
  END b5_c3_not
  PIN b5_c2
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 778.060 131.815 779.340 132.195 ;
        RECT 764.560 129.415 765.745 129.795 ;
        RECT 778.060 129.415 779.075 129.795 ;
        RECT 752.855 126.735 779.085 127.125 ;
        RECT 764.540 123.915 765.900 124.295 ;
        RECT 778.040 123.915 779.220 124.295 ;
        RECT 778.040 121.915 779.115 122.295 ;
      LAYER Metal2 ;
        RECT 765.180 129.780 765.490 129.810 ;
        RECT 765.180 123.680 765.495 129.780 ;
        RECT 778.680 121.685 779.010 132.380 ;
    END
  END b5_c2
  PIN b5_c1
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 778.000 151.620 779.280 152.000 ;
        RECT 764.500 149.220 765.685 149.600 ;
        RECT 778.000 149.220 779.015 149.600 ;
        RECT 752.795 146.540 779.025 146.930 ;
        RECT 764.480 143.720 765.840 144.100 ;
        RECT 777.980 143.720 779.160 144.100 ;
        RECT 777.980 141.720 779.055 142.100 ;
      LAYER Metal2 ;
        RECT 765.120 149.585 765.430 149.615 ;
        RECT 765.120 143.485 765.435 149.585 ;
        RECT 778.620 141.490 778.950 152.185 ;
    END
  END b5_c1
  PIN b5_c1_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 754.305 151.520 755.760 151.900 ;
        RECT 754.465 149.220 755.760 149.600 ;
        RECT 767.950 149.220 769.260 149.600 ;
        RECT 752.795 147.895 768.805 148.270 ;
        RECT 754.475 143.720 755.780 144.100 ;
        RECT 767.815 143.720 769.280 144.100 ;
        RECT 754.290 141.720 755.780 142.100 ;
      LAYER Metal2 ;
        RECT 754.595 141.010 754.950 152.095 ;
        RECT 768.105 143.440 768.435 149.635 ;
    END
  END b5_c1_not
  PIN b5_c4
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 778.020 92.320 779.300 92.700 ;
        RECT 764.520 89.920 765.705 90.300 ;
        RECT 778.020 89.920 779.035 90.300 ;
        RECT 752.815 87.240 779.045 87.630 ;
        RECT 764.500 84.420 765.860 84.800 ;
        RECT 778.000 84.420 779.180 84.800 ;
        RECT 778.000 82.420 779.075 82.800 ;
      LAYER Metal2 ;
        RECT 765.140 90.285 765.450 90.315 ;
        RECT 765.140 84.185 765.455 90.285 ;
        RECT 778.640 82.190 778.970 92.885 ;
    END
  END b5_c4
  PIN b5_p4_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.585 197.875 1143.750 198.145 ;
        RECT -21.315 109.260 -20.935 109.305 ;
        RECT -15.815 109.260 -15.435 109.305 ;
        RECT -21.365 108.945 -15.430 109.260 ;
        RECT -21.315 108.925 -20.935 108.945 ;
        RECT -15.815 108.925 -15.435 108.945 ;
        RECT -29.315 101.435 -28.225 101.815 ;
        RECT -7.815 101.770 -7.435 101.815 ;
        RECT -8.550 101.470 -7.240 101.770 ;
        RECT -7.815 101.435 -7.435 101.470 ;
        RECT -41.555 100.925 -32.095 100.935 ;
        RECT -41.555 100.585 -5.805 100.925 ;
        RECT -32.460 100.575 -5.805 100.585 ;
        RECT 174.885 89.545 175.265 89.590 ;
        RECT 180.385 89.545 180.765 89.590 ;
        RECT 567.595 89.550 567.975 89.595 ;
        RECT 573.095 89.550 573.475 89.595 ;
        RECT 763.960 89.555 764.340 89.600 ;
        RECT 769.460 89.555 769.840 89.600 ;
        RECT -71.610 89.455 -71.230 89.500 ;
        RECT -66.110 89.455 -65.730 89.500 ;
        RECT -71.660 89.140 -65.725 89.455 ;
        RECT 174.835 89.230 180.770 89.545 ;
        RECT 371.275 89.505 371.655 89.550 ;
        RECT 376.775 89.505 377.155 89.550 ;
        RECT 174.885 89.210 175.265 89.230 ;
        RECT 180.385 89.210 180.765 89.230 ;
        RECT 371.225 89.190 377.160 89.505 ;
        RECT 567.545 89.235 573.480 89.550 ;
        RECT 763.910 89.240 769.845 89.555 ;
        RECT 960.345 89.540 960.725 89.585 ;
        RECT 965.845 89.540 966.225 89.585 ;
        RECT 1156.670 89.545 1157.050 89.590 ;
        RECT 1162.170 89.545 1162.550 89.590 ;
        RECT 567.595 89.215 567.975 89.235 ;
        RECT 573.095 89.215 573.475 89.235 ;
        RECT 763.960 89.220 764.340 89.240 ;
        RECT 769.460 89.220 769.840 89.240 ;
        RECT 960.295 89.225 966.230 89.540 ;
        RECT 1156.620 89.230 1162.555 89.545 ;
        RECT 960.345 89.205 960.725 89.225 ;
        RECT 965.845 89.205 966.225 89.225 ;
        RECT 1156.670 89.210 1157.050 89.230 ;
        RECT 1162.170 89.210 1162.550 89.230 ;
        RECT 371.275 89.170 371.655 89.190 ;
        RECT 376.775 89.170 377.155 89.190 ;
        RECT -71.610 89.120 -71.230 89.140 ;
        RECT -66.110 89.120 -65.730 89.140 ;
        RECT -79.610 81.630 -78.520 82.010 ;
        RECT -58.110 81.965 -57.730 82.010 ;
        RECT -58.845 81.665 -57.535 81.965 ;
        RECT 166.885 81.720 167.975 82.100 ;
        RECT 188.385 82.055 188.765 82.100 ;
        RECT 187.650 81.755 188.960 82.055 ;
        RECT 188.385 81.720 188.765 81.755 ;
        RECT 363.275 81.680 364.365 82.060 ;
        RECT 384.775 82.015 385.155 82.060 ;
        RECT 384.040 81.715 385.350 82.015 ;
        RECT 559.595 81.725 560.685 82.105 ;
        RECT 581.095 82.060 581.475 82.105 ;
        RECT 580.360 81.760 581.670 82.060 ;
        RECT 581.095 81.725 581.475 81.760 ;
        RECT 755.960 81.730 757.050 82.110 ;
        RECT 777.460 82.065 777.840 82.110 ;
        RECT 776.725 81.765 778.035 82.065 ;
        RECT 777.460 81.730 777.840 81.765 ;
        RECT 952.345 81.715 953.435 82.095 ;
        RECT 973.845 82.050 974.225 82.095 ;
        RECT 973.110 81.750 974.420 82.050 ;
        RECT 973.845 81.715 974.225 81.750 ;
        RECT 1148.670 81.720 1149.760 82.100 ;
        RECT 1170.170 82.055 1170.550 82.100 ;
        RECT 1169.435 81.755 1170.745 82.055 ;
        RECT 1170.170 81.720 1170.550 81.755 ;
        RECT 384.775 81.680 385.155 81.715 ;
        RECT -58.110 81.630 -57.730 81.665 ;
        RECT 743.680 81.220 753.140 81.225 ;
        RECT 547.315 81.215 556.775 81.220 ;
        RECT 154.605 81.210 164.065 81.215 ;
        RECT -82.755 81.115 -56.100 81.120 ;
        RECT -91.320 80.770 -56.100 81.115 ;
        RECT 154.605 80.865 190.395 81.210 ;
        RECT 163.740 80.860 190.395 80.865 ;
        RECT 350.995 81.170 360.455 81.175 ;
        RECT 350.995 80.825 386.785 81.170 ;
        RECT 547.315 80.870 583.105 81.215 ;
        RECT 743.680 80.875 779.470 81.220 ;
        RECT 1136.390 81.210 1145.850 81.215 ;
        RECT 752.815 80.870 779.470 80.875 ;
        RECT 940.065 81.205 949.525 81.210 ;
        RECT 556.450 80.865 583.105 80.870 ;
        RECT 940.065 80.860 975.855 81.205 ;
        RECT 1136.390 80.865 1172.180 81.210 ;
        RECT 1145.525 80.860 1172.180 80.865 ;
        RECT 949.200 80.855 975.855 80.860 ;
        RECT 360.130 80.820 386.785 80.825 ;
        RECT -91.320 80.765 -82.565 80.770 ;
      LAYER Metal2 ;
        RECT -91.070 17.990 -90.775 204.535 ;
        RECT -78.995 80.770 -78.615 82.145 ;
        RECT -69.285 80.480 -68.915 89.580 ;
        RECT -58.740 80.685 -58.405 82.035 ;
        RECT -41.335 18.000 -40.985 204.525 ;
        RECT -28.700 100.575 -28.320 101.950 ;
        RECT -18.990 100.285 -18.620 109.385 ;
        RECT -8.445 100.490 -8.110 101.840 ;
        RECT 154.835 18.010 155.185 204.535 ;
        RECT 167.500 80.860 167.880 82.235 ;
        RECT 177.210 80.570 177.580 89.670 ;
        RECT 187.755 80.775 188.090 82.125 ;
        RECT 351.225 17.970 351.575 204.495 ;
        RECT 363.890 80.820 364.270 82.195 ;
        RECT 373.600 80.530 373.970 89.630 ;
        RECT 384.145 80.735 384.480 82.085 ;
        RECT 547.545 18.015 547.895 204.540 ;
        RECT 560.210 80.865 560.590 82.240 ;
        RECT 569.920 80.575 570.290 89.675 ;
        RECT 580.465 80.780 580.800 82.130 ;
        RECT 743.910 18.020 744.260 204.545 ;
        RECT 756.575 80.870 756.955 82.245 ;
        RECT 766.285 80.580 766.655 89.680 ;
        RECT 776.830 80.785 777.165 82.135 ;
        RECT 940.295 18.005 940.645 204.530 ;
        RECT 952.960 80.855 953.340 82.230 ;
        RECT 962.670 80.565 963.040 89.665 ;
        RECT 973.215 80.770 973.550 82.120 ;
        RECT 1136.620 18.010 1136.970 204.535 ;
        RECT 1149.285 80.860 1149.665 82.235 ;
        RECT 1158.995 80.570 1159.365 89.670 ;
        RECT 1169.540 80.775 1169.875 82.125 ;
    END
  END b5_p4_not
  PIN b5_p4
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.615 198.395 1143.755 198.685 ;
        RECT -42.495 113.120 -32.245 113.130 ;
        RECT -42.495 112.845 -5.805 113.120 ;
        RECT -32.460 112.835 -5.805 112.845 ;
        RECT -7.815 111.670 -7.435 111.705 ;
        RECT -29.315 111.565 -28.935 111.605 ;
        RECT -29.385 111.260 -26.550 111.565 ;
        RECT -10.570 111.360 -7.435 111.670 ;
        RECT -7.815 111.325 -7.435 111.360 ;
        RECT -29.315 111.225 -28.935 111.260 ;
        RECT -25.315 103.435 -24.225 103.815 ;
        RECT -12.770 103.435 -11.435 103.815 ;
        RECT -24.830 101.440 -11.980 101.775 ;
        RECT 742.740 93.415 752.990 93.420 ;
        RECT 546.375 93.410 556.625 93.415 ;
        RECT 153.665 93.405 163.915 93.410 ;
        RECT -82.755 93.310 -56.100 93.315 ;
        RECT -92.260 93.030 -56.100 93.310 ;
        RECT 153.665 93.125 190.395 93.405 ;
        RECT 163.740 93.120 190.395 93.125 ;
        RECT 350.055 93.365 360.305 93.370 ;
        RECT 350.055 93.085 386.785 93.365 ;
        RECT 546.375 93.130 583.105 93.410 ;
        RECT 742.740 93.135 779.470 93.415 ;
        RECT 1135.450 93.405 1145.700 93.410 ;
        RECT 752.815 93.130 779.470 93.135 ;
        RECT 939.125 93.400 949.375 93.405 ;
        RECT 556.450 93.125 583.105 93.130 ;
        RECT 939.125 93.120 975.855 93.400 ;
        RECT 1135.450 93.125 1172.180 93.405 ;
        RECT 1145.525 93.120 1172.180 93.125 ;
        RECT 949.200 93.115 975.855 93.120 ;
        RECT 360.130 93.080 386.785 93.085 ;
        RECT -92.260 93.025 -82.465 93.030 ;
        RECT 188.385 91.955 188.765 91.990 ;
        RECT 581.095 91.960 581.475 91.995 ;
        RECT 777.460 91.965 777.840 92.000 ;
        RECT -58.110 91.865 -57.730 91.900 ;
        RECT -79.610 91.760 -79.230 91.800 ;
        RECT -79.680 91.455 -76.845 91.760 ;
        RECT -60.865 91.555 -57.730 91.865 ;
        RECT 166.885 91.850 167.265 91.890 ;
        RECT -58.110 91.520 -57.730 91.555 ;
        RECT 166.815 91.545 169.650 91.850 ;
        RECT 185.630 91.645 188.765 91.955 ;
        RECT 384.775 91.915 385.155 91.950 ;
        RECT 363.275 91.810 363.655 91.850 ;
        RECT 188.385 91.610 188.765 91.645 ;
        RECT 166.885 91.510 167.265 91.545 ;
        RECT 363.205 91.505 366.040 91.810 ;
        RECT 382.020 91.605 385.155 91.915 ;
        RECT 559.595 91.855 559.975 91.895 ;
        RECT 384.775 91.570 385.155 91.605 ;
        RECT 559.525 91.550 562.360 91.855 ;
        RECT 578.340 91.650 581.475 91.960 ;
        RECT 755.960 91.860 756.340 91.900 ;
        RECT 581.095 91.615 581.475 91.650 ;
        RECT 755.890 91.555 758.725 91.860 ;
        RECT 774.705 91.655 777.840 91.965 ;
        RECT 973.845 91.950 974.225 91.985 ;
        RECT 1170.170 91.955 1170.550 91.990 ;
        RECT 952.345 91.845 952.725 91.885 ;
        RECT 777.460 91.620 777.840 91.655 ;
        RECT 559.595 91.515 559.975 91.550 ;
        RECT 755.960 91.520 756.340 91.555 ;
        RECT 952.275 91.540 955.110 91.845 ;
        RECT 971.090 91.640 974.225 91.950 ;
        RECT 1148.670 91.850 1149.050 91.890 ;
        RECT 973.845 91.605 974.225 91.640 ;
        RECT 1148.600 91.545 1151.435 91.850 ;
        RECT 1167.415 91.645 1170.550 91.955 ;
        RECT 1170.170 91.610 1170.550 91.645 ;
        RECT 952.345 91.505 952.725 91.540 ;
        RECT 1148.670 91.510 1149.050 91.545 ;
        RECT 363.275 91.470 363.655 91.505 ;
        RECT -79.610 91.420 -79.230 91.455 ;
        RECT -75.610 83.630 -74.520 84.010 ;
        RECT -63.065 83.630 -61.730 84.010 ;
        RECT 170.885 83.720 171.975 84.100 ;
        RECT 183.430 83.720 184.765 84.100 ;
        RECT 367.275 83.680 368.365 84.060 ;
        RECT 379.820 83.680 381.155 84.060 ;
        RECT 563.595 83.725 564.685 84.105 ;
        RECT 576.140 83.725 577.475 84.105 ;
        RECT 759.960 83.730 761.050 84.110 ;
        RECT 772.505 83.730 773.840 84.110 ;
        RECT 956.345 83.715 957.435 84.095 ;
        RECT 968.890 83.715 970.225 84.095 ;
        RECT 1152.670 83.720 1153.760 84.100 ;
        RECT 1165.215 83.720 1166.550 84.100 ;
        RECT -75.125 81.635 -62.275 81.970 ;
        RECT 171.370 81.725 184.220 82.060 ;
        RECT 367.760 81.685 380.610 82.020 ;
        RECT 564.080 81.730 576.930 82.065 ;
        RECT 760.445 81.735 773.295 82.070 ;
        RECT 956.830 81.720 969.680 82.055 ;
        RECT 1153.155 81.725 1166.005 82.060 ;
      LAYER Metal2 ;
        RECT -92.095 18.000 -91.755 204.535 ;
        RECT -77.210 91.335 -76.920 93.395 ;
        RECT -74.920 81.420 -74.595 84.185 ;
        RECT -68.340 81.545 -68.050 93.380 ;
        RECT -60.435 91.275 -60.125 93.790 ;
        RECT -62.985 81.420 -62.660 84.185 ;
        RECT -42.350 18.000 -41.995 204.500 ;
        RECT -26.915 111.140 -26.625 113.200 ;
        RECT -24.625 101.225 -24.300 103.990 ;
        RECT -18.045 101.350 -17.755 113.185 ;
        RECT -10.140 111.080 -9.830 113.595 ;
        RECT -12.690 101.225 -12.365 103.990 ;
        RECT 153.820 18.010 154.175 204.510 ;
        RECT 169.285 91.425 169.575 93.485 ;
        RECT 171.575 81.510 171.900 84.275 ;
        RECT 178.155 81.635 178.445 93.470 ;
        RECT 186.060 91.365 186.370 93.880 ;
        RECT 183.510 81.510 183.835 84.275 ;
        RECT 350.210 17.970 350.565 204.470 ;
        RECT 365.675 91.385 365.965 93.445 ;
        RECT 367.965 81.470 368.290 84.235 ;
        RECT 374.545 81.595 374.835 93.430 ;
        RECT 382.450 91.325 382.760 93.840 ;
        RECT 379.900 81.470 380.225 84.235 ;
        RECT 546.530 18.015 546.885 204.515 ;
        RECT 561.995 91.430 562.285 93.490 ;
        RECT 564.285 81.515 564.610 84.280 ;
        RECT 570.865 81.640 571.155 93.475 ;
        RECT 578.770 91.370 579.080 93.885 ;
        RECT 576.220 81.515 576.545 84.280 ;
        RECT 742.895 18.020 743.250 204.520 ;
        RECT 758.360 91.435 758.650 93.495 ;
        RECT 760.650 81.520 760.975 84.285 ;
        RECT 767.230 81.645 767.520 93.480 ;
        RECT 775.135 91.375 775.445 93.890 ;
        RECT 772.585 81.520 772.910 84.285 ;
        RECT 939.280 18.005 939.635 204.505 ;
        RECT 954.745 91.420 955.035 93.480 ;
        RECT 957.035 81.505 957.360 84.270 ;
        RECT 963.615 81.630 963.905 93.465 ;
        RECT 971.520 91.360 971.830 93.875 ;
        RECT 968.970 81.505 969.295 84.270 ;
        RECT 1135.605 18.010 1135.960 204.510 ;
        RECT 1151.070 91.425 1151.360 93.485 ;
        RECT 1153.360 81.510 1153.685 84.275 ;
        RECT 1159.940 81.635 1160.230 93.470 ;
        RECT 1167.845 91.365 1168.155 93.880 ;
        RECT 1165.295 81.510 1165.620 84.275 ;
    END
  END b5_p4
  PIN b5_p5_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.595 196.680 1143.745 197.005 ;
        RECT -21.285 89.535 -20.905 89.580 ;
        RECT -15.785 89.535 -15.405 89.580 ;
        RECT -21.335 89.220 -15.400 89.535 ;
        RECT -21.285 89.200 -20.905 89.220 ;
        RECT -15.785 89.200 -15.405 89.220 ;
        RECT -29.285 81.710 -28.195 82.090 ;
        RECT -7.785 82.045 -7.405 82.090 ;
        RECT -8.520 81.745 -7.210 82.045 ;
        RECT -7.785 81.710 -7.405 81.745 ;
        RECT -32.430 81.190 -5.775 81.200 ;
        RECT -39.555 80.850 -5.775 81.190 ;
        RECT -39.555 80.840 -32.270 80.850 ;
        RECT 174.815 69.715 175.195 69.760 ;
        RECT 180.315 69.715 180.695 69.760 ;
        RECT 567.525 69.720 567.905 69.765 ;
        RECT 573.025 69.720 573.405 69.765 ;
        RECT 763.890 69.725 764.270 69.770 ;
        RECT 769.390 69.725 769.770 69.770 ;
        RECT -71.680 69.625 -71.300 69.670 ;
        RECT -66.180 69.625 -65.800 69.670 ;
        RECT -71.730 69.310 -65.795 69.625 ;
        RECT 174.765 69.400 180.700 69.715 ;
        RECT 371.205 69.675 371.585 69.720 ;
        RECT 376.705 69.675 377.085 69.720 ;
        RECT 174.815 69.380 175.195 69.400 ;
        RECT 180.315 69.380 180.695 69.400 ;
        RECT 371.155 69.360 377.090 69.675 ;
        RECT 567.475 69.405 573.410 69.720 ;
        RECT 763.840 69.410 769.775 69.725 ;
        RECT 960.275 69.710 960.655 69.755 ;
        RECT 965.775 69.710 966.155 69.755 ;
        RECT 1156.600 69.715 1156.980 69.760 ;
        RECT 1162.100 69.715 1162.480 69.760 ;
        RECT 567.525 69.385 567.905 69.405 ;
        RECT 573.025 69.385 573.405 69.405 ;
        RECT 763.890 69.390 764.270 69.410 ;
        RECT 769.390 69.390 769.770 69.410 ;
        RECT 960.225 69.395 966.160 69.710 ;
        RECT 1156.550 69.400 1162.485 69.715 ;
        RECT 960.275 69.375 960.655 69.395 ;
        RECT 965.775 69.375 966.155 69.395 ;
        RECT 1156.600 69.380 1156.980 69.400 ;
        RECT 1162.100 69.380 1162.480 69.400 ;
        RECT 371.205 69.340 371.585 69.360 ;
        RECT 376.705 69.340 377.085 69.360 ;
        RECT -71.680 69.290 -71.300 69.310 ;
        RECT -66.180 69.290 -65.800 69.310 ;
        RECT -79.680 61.800 -78.590 62.180 ;
        RECT -58.180 62.135 -57.800 62.180 ;
        RECT -58.915 61.835 -57.605 62.135 ;
        RECT 166.815 61.890 167.905 62.270 ;
        RECT 188.315 62.225 188.695 62.270 ;
        RECT 187.580 61.925 188.890 62.225 ;
        RECT 188.315 61.890 188.695 61.925 ;
        RECT 363.205 61.850 364.295 62.230 ;
        RECT 384.705 62.185 385.085 62.230 ;
        RECT 383.970 61.885 385.280 62.185 ;
        RECT 559.525 61.895 560.615 62.275 ;
        RECT 581.025 62.230 581.405 62.275 ;
        RECT 580.290 61.930 581.600 62.230 ;
        RECT 581.025 61.895 581.405 61.930 ;
        RECT 755.890 61.900 756.980 62.280 ;
        RECT 777.390 62.235 777.770 62.280 ;
        RECT 776.655 61.935 777.965 62.235 ;
        RECT 777.390 61.900 777.770 61.935 ;
        RECT 952.275 61.885 953.365 62.265 ;
        RECT 973.775 62.220 974.155 62.265 ;
        RECT 973.040 61.920 974.350 62.220 ;
        RECT 973.775 61.885 974.155 61.920 ;
        RECT 1148.600 61.890 1149.690 62.270 ;
        RECT 1170.100 62.225 1170.480 62.270 ;
        RECT 1169.365 61.925 1170.675 62.225 ;
        RECT 1170.100 61.890 1170.480 61.925 ;
        RECT 384.705 61.850 385.085 61.885 ;
        RECT -58.180 61.800 -57.800 61.835 ;
        RECT 156.605 61.380 163.890 61.470 ;
        RECT -89.315 61.290 -82.585 61.305 ;
        RECT -89.315 60.955 -56.170 61.290 ;
        RECT 156.605 61.120 190.325 61.380 ;
        RECT 163.670 61.030 190.325 61.120 ;
        RECT 352.995 61.340 360.280 61.430 ;
        RECT 549.315 61.385 556.600 61.475 ;
        RECT 745.680 61.390 752.965 61.480 ;
        RECT 352.995 61.080 386.715 61.340 ;
        RECT 549.315 61.125 583.035 61.385 ;
        RECT 745.680 61.130 779.400 61.390 ;
        RECT 360.060 60.990 386.715 61.080 ;
        RECT 556.380 61.035 583.035 61.125 ;
        RECT 752.745 61.040 779.400 61.130 ;
        RECT 942.065 61.375 949.350 61.465 ;
        RECT 1138.390 61.380 1145.675 61.470 ;
        RECT 942.065 61.115 975.785 61.375 ;
        RECT 1138.390 61.120 1172.110 61.380 ;
        RECT 949.130 61.025 975.785 61.115 ;
        RECT 1145.455 61.030 1172.110 61.120 ;
        RECT -82.825 60.940 -56.170 60.955 ;
      LAYER Metal2 ;
        RECT -89.075 18.005 -88.785 204.535 ;
        RECT -79.065 60.940 -78.685 62.315 ;
        RECT -69.355 60.650 -68.985 69.750 ;
        RECT -58.810 60.855 -58.475 62.205 ;
        RECT -39.340 18.005 -38.990 204.500 ;
        RECT -28.670 80.850 -28.290 82.225 ;
        RECT -18.960 80.560 -18.590 89.660 ;
        RECT -8.415 80.765 -8.080 82.115 ;
        RECT 156.830 18.015 157.180 204.510 ;
        RECT 167.430 61.030 167.810 62.405 ;
        RECT 177.140 60.740 177.510 69.840 ;
        RECT 187.685 60.945 188.020 62.295 ;
        RECT 353.220 17.975 353.570 204.470 ;
        RECT 363.820 60.990 364.200 62.365 ;
        RECT 373.530 60.700 373.900 69.800 ;
        RECT 384.075 60.905 384.410 62.255 ;
        RECT 549.540 18.020 549.890 204.515 ;
        RECT 560.140 61.035 560.520 62.410 ;
        RECT 569.850 60.745 570.220 69.845 ;
        RECT 580.395 60.950 580.730 62.300 ;
        RECT 745.905 18.025 746.255 204.520 ;
        RECT 756.505 61.040 756.885 62.415 ;
        RECT 766.215 60.750 766.585 69.850 ;
        RECT 776.760 60.955 777.095 62.305 ;
        RECT 942.290 18.010 942.640 204.505 ;
        RECT 952.890 61.025 953.270 62.400 ;
        RECT 962.600 60.735 962.970 69.835 ;
        RECT 973.145 60.940 973.480 62.290 ;
        RECT 1138.615 18.015 1138.965 204.510 ;
        RECT 1149.215 61.030 1149.595 62.405 ;
        RECT 1158.925 60.740 1159.295 69.840 ;
        RECT 1169.470 60.945 1169.805 62.295 ;
    END
  END b5_p5_not
  PIN b5_c5_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 754.255 72.390 755.710 72.770 ;
        RECT 754.415 70.090 755.710 70.470 ;
        RECT 767.900 70.090 769.210 70.470 ;
        RECT 752.745 68.765 768.755 69.140 ;
        RECT 754.425 64.590 755.730 64.970 ;
        RECT 767.765 64.590 769.230 64.970 ;
        RECT 754.240 62.590 755.730 62.970 ;
      LAYER Metal2 ;
        RECT 754.545 61.880 754.900 72.965 ;
        RECT 768.055 64.310 768.385 70.505 ;
    END
  END b5_c5_not
  PIN b5_c5
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 777.950 72.490 779.230 72.870 ;
        RECT 764.450 70.090 765.635 70.470 ;
        RECT 777.950 70.090 778.965 70.470 ;
        RECT 752.745 67.410 778.975 67.800 ;
        RECT 764.430 64.590 765.790 64.970 ;
        RECT 777.930 64.590 779.110 64.970 ;
        RECT 777.930 62.590 779.005 62.970 ;
      LAYER Metal2 ;
        RECT 765.070 70.455 765.380 70.485 ;
        RECT 765.070 64.355 765.385 70.455 ;
        RECT 778.570 62.360 778.900 73.055 ;
    END
  END b5_c5
  PIN b5_c6_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 754.325 52.670 755.780 53.050 ;
        RECT 754.485 50.370 755.780 50.750 ;
        RECT 767.970 50.370 769.280 50.750 ;
        RECT 752.815 49.045 768.825 49.420 ;
        RECT 754.495 44.870 755.800 45.250 ;
        RECT 767.835 44.870 769.300 45.250 ;
        RECT 754.310 42.870 755.800 43.250 ;
      LAYER Metal2 ;
        RECT 754.615 42.160 754.970 53.245 ;
        RECT 768.125 44.590 768.455 50.785 ;
    END
  END b5_c6_not
  PIN b5_c6
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 778.020 52.770 779.300 53.150 ;
        RECT 764.520 50.370 765.705 50.750 ;
        RECT 778.020 50.370 779.035 50.750 ;
        RECT 752.815 47.690 779.045 48.080 ;
        RECT 764.500 44.870 765.860 45.250 ;
        RECT 778.000 44.870 779.180 45.250 ;
        RECT 778.000 42.870 779.075 43.250 ;
      LAYER Metal2 ;
        RECT 765.140 50.735 765.450 50.765 ;
        RECT 765.140 44.635 765.455 50.735 ;
        RECT 778.640 42.640 778.970 53.335 ;
    END
  END b5_c6
  PIN vss
    ANTENNADIFFAREA 0.514800 ;
    PORT
      LAYER Pwell ;
        RECT 664.010 0.270 679.470 7.970 ;
      LAYER Metal1 ;
        RECT 664.010 1.165 667.675 1.175 ;
        RECT 678.290 1.170 678.670 7.000 ;
        RECT 677.920 1.165 679.040 1.170 ;
        RECT 664.010 0.270 679.040 1.165 ;
    END
    PORT
      LAYER Pwell ;
        RECT 1056.690 0.270 1072.150 7.970 ;
      LAYER Metal1 ;
        RECT 1056.690 1.165 1060.355 1.175 ;
        RECT 1070.970 1.170 1071.350 7.000 ;
        RECT 1070.600 1.165 1071.720 1.170 ;
        RECT 1056.690 0.270 1071.720 1.165 ;
    END
    PORT
      LAYER Pwell ;
        RECT 1253.030 0.270 1268.490 7.970 ;
      LAYER Metal1 ;
        RECT 1253.030 1.165 1256.695 1.175 ;
        RECT 1267.310 1.170 1267.690 7.000 ;
        RECT 1266.940 1.165 1268.060 1.170 ;
        RECT 1253.030 0.270 1268.060 1.165 ;
    END
    PORT
      LAYER Pwell ;
        RECT 74.870 0.285 90.330 7.985 ;
      LAYER Metal1 ;
        RECT 74.870 1.180 78.535 1.190 ;
        RECT 89.150 1.185 89.530 7.015 ;
        RECT 88.780 1.180 89.900 1.185 ;
        RECT 74.870 0.285 89.900 1.180 ;
    END
    PORT
      LAYER Pwell ;
        RECT 271.235 0.285 286.695 7.985 ;
      LAYER Metal1 ;
        RECT 271.235 1.180 274.900 1.190 ;
        RECT 285.515 1.185 285.895 7.015 ;
        RECT 285.145 1.180 286.265 1.185 ;
        RECT 271.235 0.285 286.265 1.180 ;
    END
    PORT
      LAYER Pwell ;
        RECT 467.635 0.235 483.095 7.935 ;
      LAYER Metal1 ;
        RECT 467.635 1.130 471.300 1.140 ;
        RECT 481.915 1.135 482.295 6.965 ;
        RECT 481.545 1.130 482.665 1.135 ;
        RECT 467.635 0.235 482.665 1.130 ;
    END
    PORT
      LAYER Pwell ;
        RECT 860.350 0.270 875.810 7.970 ;
      LAYER Metal1 ;
        RECT 860.350 1.165 864.015 1.175 ;
        RECT 874.630 1.170 875.010 7.000 ;
        RECT 874.260 1.165 875.380 1.170 ;
        RECT 860.350 0.270 875.380 1.165 ;
    END
  END vss
  PIN vdd
    ANTENNADIFFAREA 0.514800 ;
    PORT
      LAYER Nwell ;
        RECT 664.010 7.970 679.470 16.195 ;
      LAYER Metal1 ;
        RECT 664.010 15.295 679.040 16.195 ;
        RECT 678.290 8.135 678.670 15.295 ;
    END
    PORT
      LAYER Nwell ;
        RECT 860.350 7.970 875.810 16.195 ;
      LAYER Metal1 ;
        RECT 860.350 15.295 875.380 16.195 ;
        RECT 874.630 8.135 875.010 15.295 ;
    END
    PORT
      LAYER Nwell ;
        RECT 1056.690 7.970 1072.150 16.195 ;
      LAYER Metal1 ;
        RECT 1056.690 15.295 1071.720 16.195 ;
        RECT 1070.970 8.135 1071.350 15.295 ;
    END
    PORT
      LAYER Nwell ;
        RECT 1253.030 7.970 1268.490 16.195 ;
      LAYER Metal1 ;
        RECT 1253.030 15.295 1268.060 16.195 ;
        RECT 1267.310 8.135 1267.690 15.295 ;
    END
    PORT
      LAYER Nwell ;
        RECT 74.870 7.985 90.330 16.210 ;
      LAYER Metal1 ;
        RECT 74.870 15.310 89.900 16.210 ;
        RECT 89.150 8.150 89.530 15.310 ;
    END
    PORT
      LAYER Nwell ;
        RECT 271.235 7.985 286.695 16.210 ;
      LAYER Metal1 ;
        RECT 271.235 15.310 286.265 16.210 ;
        RECT 285.515 8.150 285.895 15.310 ;
    END
    PORT
      LAYER Nwell ;
        RECT 467.635 7.935 483.095 16.160 ;
      LAYER Metal1 ;
        RECT 467.635 15.260 482.665 16.160 ;
        RECT 481.915 8.100 482.295 15.260 ;
    END
  END vdd
  PIN b5_p3_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.660 198.985 1143.755 199.315 ;
        RECT -21.245 129.030 -20.865 129.075 ;
        RECT -15.745 129.030 -15.365 129.075 ;
        RECT -21.295 128.715 -15.360 129.030 ;
        RECT -21.245 128.695 -20.865 128.715 ;
        RECT -15.745 128.695 -15.365 128.715 ;
        RECT -29.245 121.205 -28.155 121.585 ;
        RECT -7.745 121.540 -7.365 121.585 ;
        RECT -8.480 121.240 -7.170 121.540 ;
        RECT -7.745 121.205 -7.365 121.240 ;
        RECT -32.390 120.670 -5.735 120.695 ;
        RECT -43.560 120.345 -5.735 120.670 ;
        RECT -43.560 120.320 -32.085 120.345 ;
        RECT 174.855 109.270 175.235 109.315 ;
        RECT 180.355 109.270 180.735 109.315 ;
        RECT 567.565 109.275 567.945 109.320 ;
        RECT 573.065 109.275 573.445 109.320 ;
        RECT 763.930 109.280 764.310 109.325 ;
        RECT 769.430 109.280 769.810 109.325 ;
        RECT -71.640 109.180 -71.260 109.225 ;
        RECT -66.140 109.180 -65.760 109.225 ;
        RECT -71.690 108.865 -65.755 109.180 ;
        RECT 174.805 108.955 180.740 109.270 ;
        RECT 371.245 109.230 371.625 109.275 ;
        RECT 376.745 109.230 377.125 109.275 ;
        RECT 174.855 108.935 175.235 108.955 ;
        RECT 180.355 108.935 180.735 108.955 ;
        RECT 371.195 108.915 377.130 109.230 ;
        RECT 567.515 108.960 573.450 109.275 ;
        RECT 763.880 108.965 769.815 109.280 ;
        RECT 960.315 109.265 960.695 109.310 ;
        RECT 965.815 109.265 966.195 109.310 ;
        RECT 1156.640 109.270 1157.020 109.315 ;
        RECT 1162.140 109.270 1162.520 109.315 ;
        RECT 567.565 108.940 567.945 108.960 ;
        RECT 573.065 108.940 573.445 108.960 ;
        RECT 763.930 108.945 764.310 108.965 ;
        RECT 769.430 108.945 769.810 108.965 ;
        RECT 960.265 108.950 966.200 109.265 ;
        RECT 1156.590 108.955 1162.525 109.270 ;
        RECT 960.315 108.930 960.695 108.950 ;
        RECT 965.815 108.930 966.195 108.950 ;
        RECT 1156.640 108.935 1157.020 108.955 ;
        RECT 1162.140 108.935 1162.520 108.955 ;
        RECT 371.245 108.895 371.625 108.915 ;
        RECT 376.745 108.895 377.125 108.915 ;
        RECT -71.640 108.845 -71.260 108.865 ;
        RECT -66.140 108.845 -65.760 108.865 ;
        RECT -79.640 101.355 -78.550 101.735 ;
        RECT -58.140 101.690 -57.760 101.735 ;
        RECT -58.875 101.390 -57.565 101.690 ;
        RECT 166.855 101.445 167.945 101.825 ;
        RECT 188.355 101.780 188.735 101.825 ;
        RECT 187.620 101.480 188.930 101.780 ;
        RECT 188.355 101.445 188.735 101.480 ;
        RECT 363.245 101.405 364.335 101.785 ;
        RECT 384.745 101.740 385.125 101.785 ;
        RECT 384.010 101.440 385.320 101.740 ;
        RECT 559.565 101.450 560.655 101.830 ;
        RECT 581.065 101.785 581.445 101.830 ;
        RECT 580.330 101.485 581.640 101.785 ;
        RECT 581.065 101.450 581.445 101.485 ;
        RECT 755.930 101.455 757.020 101.835 ;
        RECT 777.430 101.790 777.810 101.835 ;
        RECT 776.695 101.490 778.005 101.790 ;
        RECT 777.430 101.455 777.810 101.490 ;
        RECT 952.315 101.440 953.405 101.820 ;
        RECT 973.815 101.775 974.195 101.820 ;
        RECT 973.080 101.475 974.390 101.775 ;
        RECT 973.815 101.440 974.195 101.475 ;
        RECT 1148.640 101.445 1149.730 101.825 ;
        RECT 1170.140 101.780 1170.520 101.825 ;
        RECT 1169.405 101.480 1170.715 101.780 ;
        RECT 1170.140 101.445 1170.520 101.480 ;
        RECT 384.745 101.405 385.125 101.440 ;
        RECT -58.140 101.355 -57.760 101.390 ;
        RECT 152.600 100.935 164.075 100.950 ;
        RECT 545.310 100.940 556.785 100.955 ;
        RECT 741.675 100.945 753.150 100.960 ;
        RECT -93.325 100.845 -82.550 100.850 ;
        RECT -93.325 100.500 -56.130 100.845 ;
        RECT 152.600 100.600 190.365 100.935 ;
        RECT 163.710 100.585 190.365 100.600 ;
        RECT 348.990 100.895 360.465 100.910 ;
        RECT 348.990 100.560 386.755 100.895 ;
        RECT 545.310 100.605 583.075 100.940 ;
        RECT 741.675 100.610 779.440 100.945 ;
        RECT 556.420 100.590 583.075 100.605 ;
        RECT 752.785 100.595 779.440 100.610 ;
        RECT 938.060 100.930 949.535 100.945 ;
        RECT 1134.385 100.935 1145.860 100.950 ;
        RECT 938.060 100.595 975.825 100.930 ;
        RECT 1134.385 100.600 1172.150 100.935 ;
        RECT 949.170 100.580 975.825 100.595 ;
        RECT 1145.495 100.585 1172.150 100.600 ;
        RECT 360.100 100.545 386.755 100.560 ;
        RECT -82.785 100.495 -56.130 100.500 ;
      LAYER Metal2 ;
        RECT -93.200 17.985 -92.805 204.520 ;
        RECT -79.025 100.495 -78.645 101.870 ;
        RECT -69.315 100.205 -68.945 109.305 ;
        RECT -58.770 100.410 -58.435 101.760 ;
        RECT -43.415 18.010 -43.095 204.525 ;
        RECT -28.630 120.345 -28.250 121.720 ;
        RECT -18.920 120.055 -18.550 129.155 ;
        RECT -8.375 120.260 -8.040 121.610 ;
        RECT 152.755 18.020 153.075 204.535 ;
        RECT 167.470 100.585 167.850 101.960 ;
        RECT 177.180 100.295 177.550 109.395 ;
        RECT 187.725 100.500 188.060 101.850 ;
        RECT 349.145 17.980 349.465 204.495 ;
        RECT 363.860 100.545 364.240 101.920 ;
        RECT 373.570 100.255 373.940 109.355 ;
        RECT 384.115 100.460 384.450 101.810 ;
        RECT 545.465 18.025 545.785 204.540 ;
        RECT 560.180 100.590 560.560 101.965 ;
        RECT 569.890 100.300 570.260 109.400 ;
        RECT 580.435 100.505 580.770 101.855 ;
        RECT 741.830 18.030 742.150 204.545 ;
        RECT 756.545 100.595 756.925 101.970 ;
        RECT 766.255 100.305 766.625 109.405 ;
        RECT 776.800 100.510 777.135 101.860 ;
        RECT 938.215 18.015 938.535 204.530 ;
        RECT 952.930 100.580 953.310 101.955 ;
        RECT 962.640 100.290 963.010 109.390 ;
        RECT 973.185 100.495 973.520 101.845 ;
        RECT 1134.540 18.020 1134.860 204.535 ;
        RECT 1149.255 100.585 1149.635 101.960 ;
        RECT 1158.965 100.295 1159.335 109.395 ;
        RECT 1169.510 100.500 1169.845 101.850 ;
    END
  END b5_p3_not
  PIN b5_p5
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.570 197.315 1143.755 197.590 ;
        RECT -32.430 93.320 -5.775 93.395 ;
        RECT -40.525 93.110 -5.775 93.320 ;
        RECT -40.525 93.035 -32.320 93.110 ;
        RECT -7.785 91.945 -7.405 91.980 ;
        RECT -29.285 91.840 -28.905 91.880 ;
        RECT -29.355 91.535 -26.520 91.840 ;
        RECT -10.540 91.635 -7.405 91.945 ;
        RECT -7.785 91.600 -7.405 91.635 ;
        RECT -29.285 91.500 -28.905 91.535 ;
        RECT -25.285 83.710 -24.195 84.090 ;
        RECT -12.740 83.710 -11.405 84.090 ;
        RECT -24.800 81.715 -11.950 82.050 ;
        RECT 155.635 73.575 163.840 73.600 ;
        RECT 548.345 73.580 556.550 73.605 ;
        RECT 744.710 73.585 752.915 73.610 ;
        RECT -90.290 73.485 -82.485 73.500 ;
        RECT -90.290 73.215 -56.170 73.485 ;
        RECT 155.635 73.315 190.325 73.575 ;
        RECT 163.670 73.290 190.325 73.315 ;
        RECT 352.025 73.535 360.230 73.560 ;
        RECT 352.025 73.275 386.715 73.535 ;
        RECT 548.345 73.320 583.035 73.580 ;
        RECT 744.710 73.325 779.400 73.585 ;
        RECT 556.380 73.295 583.035 73.320 ;
        RECT 752.745 73.300 779.400 73.325 ;
        RECT 941.095 73.570 949.300 73.595 ;
        RECT 1137.420 73.575 1145.625 73.600 ;
        RECT 941.095 73.310 975.785 73.570 ;
        RECT 1137.420 73.315 1172.110 73.575 ;
        RECT 949.130 73.285 975.785 73.310 ;
        RECT 1145.455 73.290 1172.110 73.315 ;
        RECT 360.060 73.250 386.715 73.275 ;
        RECT -82.825 73.200 -56.170 73.215 ;
        RECT 188.315 72.125 188.695 72.160 ;
        RECT 581.025 72.130 581.405 72.165 ;
        RECT 777.390 72.135 777.770 72.170 ;
        RECT -58.180 72.035 -57.800 72.070 ;
        RECT -79.680 71.930 -79.300 71.970 ;
        RECT -79.750 71.625 -76.915 71.930 ;
        RECT -60.935 71.725 -57.800 72.035 ;
        RECT 166.815 72.020 167.195 72.060 ;
        RECT -58.180 71.690 -57.800 71.725 ;
        RECT 166.745 71.715 169.580 72.020 ;
        RECT 185.560 71.815 188.695 72.125 ;
        RECT 384.705 72.085 385.085 72.120 ;
        RECT 363.205 71.980 363.585 72.020 ;
        RECT 188.315 71.780 188.695 71.815 ;
        RECT 166.815 71.680 167.195 71.715 ;
        RECT 363.135 71.675 365.970 71.980 ;
        RECT 381.950 71.775 385.085 72.085 ;
        RECT 559.525 72.025 559.905 72.065 ;
        RECT 384.705 71.740 385.085 71.775 ;
        RECT 559.455 71.720 562.290 72.025 ;
        RECT 578.270 71.820 581.405 72.130 ;
        RECT 755.890 72.030 756.270 72.070 ;
        RECT 581.025 71.785 581.405 71.820 ;
        RECT 755.820 71.725 758.655 72.030 ;
        RECT 774.635 71.825 777.770 72.135 ;
        RECT 973.775 72.120 974.155 72.155 ;
        RECT 1170.100 72.125 1170.480 72.160 ;
        RECT 952.275 72.015 952.655 72.055 ;
        RECT 777.390 71.790 777.770 71.825 ;
        RECT 559.525 71.685 559.905 71.720 ;
        RECT 755.890 71.690 756.270 71.725 ;
        RECT 952.205 71.710 955.040 72.015 ;
        RECT 971.020 71.810 974.155 72.120 ;
        RECT 1148.600 72.020 1148.980 72.060 ;
        RECT 973.775 71.775 974.155 71.810 ;
        RECT 1148.530 71.715 1151.365 72.020 ;
        RECT 1167.345 71.815 1170.480 72.125 ;
        RECT 1170.100 71.780 1170.480 71.815 ;
        RECT 952.275 71.675 952.655 71.710 ;
        RECT 1148.600 71.680 1148.980 71.715 ;
        RECT 363.205 71.640 363.585 71.675 ;
        RECT -79.680 71.590 -79.300 71.625 ;
        RECT -75.680 63.800 -74.590 64.180 ;
        RECT -63.135 63.800 -61.800 64.180 ;
        RECT 170.815 63.890 171.905 64.270 ;
        RECT 183.360 63.890 184.695 64.270 ;
        RECT 367.205 63.850 368.295 64.230 ;
        RECT 379.750 63.850 381.085 64.230 ;
        RECT 563.525 63.895 564.615 64.275 ;
        RECT 576.070 63.895 577.405 64.275 ;
        RECT 759.890 63.900 760.980 64.280 ;
        RECT 772.435 63.900 773.770 64.280 ;
        RECT 956.275 63.885 957.365 64.265 ;
        RECT 968.820 63.885 970.155 64.265 ;
        RECT 1152.600 63.890 1153.690 64.270 ;
        RECT 1165.145 63.890 1166.480 64.270 ;
        RECT -75.195 61.805 -62.345 62.140 ;
        RECT 171.300 61.895 184.150 62.230 ;
        RECT 367.690 61.855 380.540 62.190 ;
        RECT 564.010 61.900 576.860 62.235 ;
        RECT 760.375 61.905 773.225 62.240 ;
        RECT 956.760 61.890 969.610 62.225 ;
        RECT 1153.085 61.895 1165.935 62.230 ;
      LAYER Metal2 ;
        RECT -90.060 18.000 -89.775 204.530 ;
        RECT -77.280 71.505 -76.990 73.565 ;
        RECT -74.990 61.590 -74.665 64.355 ;
        RECT -68.410 61.715 -68.120 73.550 ;
        RECT -60.505 71.445 -60.195 73.960 ;
        RECT -63.055 61.590 -62.730 64.355 ;
        RECT -40.320 18.000 -39.995 204.490 ;
        RECT -26.885 91.415 -26.595 93.475 ;
        RECT -24.595 81.500 -24.270 84.265 ;
        RECT -18.015 81.625 -17.725 93.460 ;
        RECT -10.110 91.355 -9.800 93.870 ;
        RECT -12.660 81.500 -12.335 84.265 ;
        RECT 155.850 18.010 156.175 204.500 ;
        RECT 169.215 71.595 169.505 73.655 ;
        RECT 171.505 61.680 171.830 64.445 ;
        RECT 178.085 61.805 178.375 73.640 ;
        RECT 185.990 71.535 186.300 74.050 ;
        RECT 183.440 61.680 183.765 64.445 ;
        RECT 352.240 17.970 352.565 204.460 ;
        RECT 365.605 71.555 365.895 73.615 ;
        RECT 367.895 61.640 368.220 64.405 ;
        RECT 374.475 61.765 374.765 73.600 ;
        RECT 382.380 71.495 382.690 74.010 ;
        RECT 379.830 61.640 380.155 64.405 ;
        RECT 548.560 18.015 548.885 204.505 ;
        RECT 561.925 71.600 562.215 73.660 ;
        RECT 564.215 61.685 564.540 64.450 ;
        RECT 570.795 61.810 571.085 73.645 ;
        RECT 578.700 71.540 579.010 74.055 ;
        RECT 576.150 61.685 576.475 64.450 ;
        RECT 744.925 18.020 745.250 204.510 ;
        RECT 758.290 71.605 758.580 73.665 ;
        RECT 760.580 61.690 760.905 64.455 ;
        RECT 767.160 61.815 767.450 73.650 ;
        RECT 775.065 71.545 775.375 74.060 ;
        RECT 772.515 61.690 772.840 64.455 ;
        RECT 941.310 18.005 941.635 204.495 ;
        RECT 954.675 71.590 954.965 73.650 ;
        RECT 956.965 61.675 957.290 64.440 ;
        RECT 963.545 61.800 963.835 73.635 ;
        RECT 971.450 71.530 971.760 74.045 ;
        RECT 968.900 61.675 969.225 64.440 ;
        RECT 1137.635 18.010 1137.960 204.500 ;
        RECT 1151.000 71.595 1151.290 73.655 ;
        RECT 1153.290 61.680 1153.615 64.445 ;
        RECT 1159.870 61.805 1160.160 73.640 ;
        RECT 1167.775 71.535 1168.085 74.050 ;
        RECT 1165.225 61.680 1165.550 64.445 ;
    END
  END b5_p5
  PIN b5_p6_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.585 195.625 1143.760 195.895 ;
        RECT -21.355 69.705 -20.975 69.750 ;
        RECT -15.855 69.705 -15.475 69.750 ;
        RECT -21.405 69.390 -15.470 69.705 ;
        RECT -21.355 69.370 -20.975 69.390 ;
        RECT -15.855 69.370 -15.475 69.390 ;
        RECT -29.355 61.880 -28.265 62.260 ;
        RECT -7.855 62.215 -7.475 62.260 ;
        RECT -8.590 61.915 -7.280 62.215 ;
        RECT -7.855 61.880 -7.475 61.915 ;
        RECT -37.535 61.370 -31.845 61.390 ;
        RECT -37.535 61.040 -5.845 61.370 ;
        RECT -32.500 61.020 -5.845 61.040 ;
        RECT 174.885 49.995 175.265 50.040 ;
        RECT 180.385 49.995 180.765 50.040 ;
        RECT 567.595 50.000 567.975 50.045 ;
        RECT 573.095 50.000 573.475 50.045 ;
        RECT 763.960 50.005 764.340 50.050 ;
        RECT 769.460 50.005 769.840 50.050 ;
        RECT -71.610 49.905 -71.230 49.950 ;
        RECT -66.110 49.905 -65.730 49.950 ;
        RECT -71.660 49.590 -65.725 49.905 ;
        RECT 174.835 49.680 180.770 49.995 ;
        RECT 371.275 49.955 371.655 50.000 ;
        RECT 376.775 49.955 377.155 50.000 ;
        RECT 174.885 49.660 175.265 49.680 ;
        RECT 180.385 49.660 180.765 49.680 ;
        RECT 371.225 49.640 377.160 49.955 ;
        RECT 567.545 49.685 573.480 50.000 ;
        RECT 763.910 49.690 769.845 50.005 ;
        RECT 960.345 49.990 960.725 50.035 ;
        RECT 965.845 49.990 966.225 50.035 ;
        RECT 1156.670 49.995 1157.050 50.040 ;
        RECT 1162.170 49.995 1162.550 50.040 ;
        RECT 567.595 49.665 567.975 49.685 ;
        RECT 573.095 49.665 573.475 49.685 ;
        RECT 763.960 49.670 764.340 49.690 ;
        RECT 769.460 49.670 769.840 49.690 ;
        RECT 960.295 49.675 966.230 49.990 ;
        RECT 1156.620 49.680 1162.555 49.995 ;
        RECT 960.345 49.655 960.725 49.675 ;
        RECT 965.845 49.655 966.225 49.675 ;
        RECT 1156.670 49.660 1157.050 49.680 ;
        RECT 1162.170 49.660 1162.550 49.680 ;
        RECT 371.275 49.620 371.655 49.640 ;
        RECT 376.775 49.620 377.155 49.640 ;
        RECT -71.610 49.570 -71.230 49.590 ;
        RECT -66.110 49.570 -65.730 49.590 ;
        RECT -79.610 42.080 -78.520 42.460 ;
        RECT -58.110 42.415 -57.730 42.460 ;
        RECT -58.845 42.115 -57.535 42.415 ;
        RECT 166.885 42.170 167.975 42.550 ;
        RECT 188.385 42.505 188.765 42.550 ;
        RECT 187.650 42.205 188.960 42.505 ;
        RECT 188.385 42.170 188.765 42.205 ;
        RECT 363.275 42.130 364.365 42.510 ;
        RECT 384.775 42.465 385.155 42.510 ;
        RECT 384.040 42.165 385.350 42.465 ;
        RECT 559.595 42.175 560.685 42.555 ;
        RECT 581.095 42.510 581.475 42.555 ;
        RECT 580.360 42.210 581.670 42.510 ;
        RECT 581.095 42.175 581.475 42.210 ;
        RECT 755.960 42.180 757.050 42.560 ;
        RECT 777.460 42.515 777.840 42.560 ;
        RECT 776.725 42.215 778.035 42.515 ;
        RECT 777.460 42.180 777.840 42.215 ;
        RECT 952.345 42.165 953.435 42.545 ;
        RECT 973.845 42.500 974.225 42.545 ;
        RECT 973.110 42.200 974.420 42.500 ;
        RECT 973.845 42.165 974.225 42.200 ;
        RECT 1148.670 42.170 1149.760 42.550 ;
        RECT 1170.170 42.505 1170.550 42.550 ;
        RECT 1169.435 42.205 1170.745 42.505 ;
        RECT 1170.170 42.170 1170.550 42.205 ;
        RECT 384.775 42.130 385.155 42.165 ;
        RECT -58.110 42.080 -57.730 42.115 ;
        RECT 158.625 41.660 164.315 41.670 ;
        RECT 551.335 41.665 557.025 41.675 ;
        RECT 747.700 41.670 753.390 41.680 ;
        RECT -87.300 41.220 -56.100 41.570 ;
        RECT 158.625 41.320 190.395 41.660 ;
        RECT 163.740 41.310 190.395 41.320 ;
        RECT 355.015 41.620 360.705 41.630 ;
        RECT 355.015 41.280 386.785 41.620 ;
        RECT 551.335 41.325 583.105 41.665 ;
        RECT 747.700 41.330 779.470 41.670 ;
        RECT 556.450 41.315 583.105 41.325 ;
        RECT 752.815 41.320 779.470 41.330 ;
        RECT 944.085 41.655 949.775 41.665 ;
        RECT 1140.410 41.660 1146.100 41.670 ;
        RECT 944.085 41.315 975.855 41.655 ;
        RECT 1140.410 41.320 1172.180 41.660 ;
        RECT 949.200 41.305 975.855 41.315 ;
        RECT 1145.525 41.310 1172.180 41.320 ;
        RECT 360.130 41.270 386.785 41.280 ;
      LAYER Metal2 ;
        RECT -87.120 18.000 -86.795 204.530 ;
        RECT -78.995 41.220 -78.615 42.595 ;
        RECT -69.285 40.930 -68.915 50.030 ;
        RECT -58.740 41.135 -58.405 42.485 ;
        RECT -37.370 18.000 -37.040 204.525 ;
        RECT -28.740 61.020 -28.360 62.395 ;
        RECT -19.030 60.730 -18.660 69.830 ;
        RECT -8.485 60.935 -8.150 62.285 ;
        RECT 158.800 18.010 159.130 204.535 ;
        RECT 167.500 41.310 167.880 42.685 ;
        RECT 177.210 41.020 177.580 50.120 ;
        RECT 187.755 41.225 188.090 42.575 ;
        RECT 355.190 17.970 355.520 204.495 ;
        RECT 363.890 41.270 364.270 42.645 ;
        RECT 373.600 40.980 373.970 50.080 ;
        RECT 384.145 41.185 384.480 42.535 ;
        RECT 551.510 18.015 551.840 204.540 ;
        RECT 560.210 41.315 560.590 42.690 ;
        RECT 569.920 41.025 570.290 50.125 ;
        RECT 580.465 41.230 580.800 42.580 ;
        RECT 747.875 18.020 748.205 204.545 ;
        RECT 756.575 41.320 756.955 42.695 ;
        RECT 766.285 41.030 766.655 50.130 ;
        RECT 776.830 41.235 777.165 42.585 ;
        RECT 944.260 18.005 944.590 204.530 ;
        RECT 952.960 41.305 953.340 42.680 ;
        RECT 962.670 41.015 963.040 50.115 ;
        RECT 973.215 41.220 973.550 42.570 ;
        RECT 1140.585 18.010 1140.915 204.535 ;
        RECT 1149.285 41.310 1149.665 42.685 ;
        RECT 1158.995 41.020 1159.365 50.120 ;
        RECT 1169.540 41.225 1169.875 42.575 ;
    END
  END b5_p6_not
  PIN b6_c4_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 950.710 92.205 952.165 92.585 ;
        RECT 950.870 89.905 952.165 90.285 ;
        RECT 964.355 89.905 965.665 90.285 ;
        RECT 949.200 88.580 965.210 88.955 ;
        RECT 950.880 84.405 952.185 84.785 ;
        RECT 964.220 84.405 965.685 84.785 ;
        RECT 950.695 82.405 952.185 82.785 ;
      LAYER Metal2 ;
        RECT 951.000 81.695 951.355 92.780 ;
        RECT 964.510 84.125 964.840 90.320 ;
    END
  END b6_c4_not
  PIN b6_c4
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 974.405 92.305 975.685 92.685 ;
        RECT 960.905 89.905 962.090 90.285 ;
        RECT 974.405 89.905 975.420 90.285 ;
        RECT 949.200 87.225 975.430 87.615 ;
        RECT 960.885 84.405 962.245 84.785 ;
        RECT 974.385 84.405 975.565 84.785 ;
        RECT 974.385 82.405 975.460 82.785 ;
      LAYER Metal2 ;
        RECT 961.525 90.270 961.835 90.300 ;
        RECT 961.525 84.170 961.840 90.270 ;
        RECT 975.025 82.175 975.355 92.870 ;
    END
  END b6_c4
  PIN b6_c5_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 950.640 72.375 952.095 72.755 ;
        RECT 950.800 70.075 952.095 70.455 ;
        RECT 964.285 70.075 965.595 70.455 ;
        RECT 949.130 68.750 965.140 69.125 ;
        RECT 950.810 64.575 952.115 64.955 ;
        RECT 964.150 64.575 965.615 64.955 ;
        RECT 950.625 62.575 952.115 62.955 ;
      LAYER Metal2 ;
        RECT 950.930 61.865 951.285 72.950 ;
        RECT 964.440 64.295 964.770 70.490 ;
    END
  END b6_c5_not
  PIN b6_c5
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 974.335 72.475 975.615 72.855 ;
        RECT 960.835 70.075 962.020 70.455 ;
        RECT 974.335 70.075 975.350 70.455 ;
        RECT 949.130 67.395 975.360 67.785 ;
        RECT 960.815 64.575 962.175 64.955 ;
        RECT 974.315 64.575 975.495 64.955 ;
        RECT 974.315 62.575 975.390 62.955 ;
      LAYER Metal2 ;
        RECT 961.455 70.440 961.765 70.470 ;
        RECT 961.455 64.340 961.770 70.440 ;
        RECT 974.955 62.345 975.285 73.040 ;
    END
  END b6_c5
  PIN b6_c6_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 950.710 52.655 952.165 53.035 ;
        RECT 950.870 50.355 952.165 50.735 ;
        RECT 964.355 50.355 965.665 50.735 ;
        RECT 949.200 49.030 965.210 49.405 ;
        RECT 950.880 44.855 952.185 45.235 ;
        RECT 964.220 44.855 965.685 45.235 ;
        RECT 950.695 42.855 952.185 43.235 ;
      LAYER Metal2 ;
        RECT 951.000 42.145 951.355 53.230 ;
        RECT 964.510 44.575 964.840 50.770 ;
    END
  END b6_c6_not
  PIN b6_c6
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 974.405 52.755 975.685 53.135 ;
        RECT 960.905 50.355 962.090 50.735 ;
        RECT 974.405 50.355 975.420 50.735 ;
        RECT 949.200 47.675 975.430 48.065 ;
        RECT 960.885 44.855 962.245 45.235 ;
        RECT 974.385 44.855 975.565 45.235 ;
        RECT 974.385 42.855 975.460 43.235 ;
      LAYER Metal2 ;
        RECT 961.525 50.720 961.835 50.750 ;
        RECT 961.525 44.620 961.840 50.720 ;
        RECT 975.025 42.625 975.355 53.320 ;
    END
  END b6_c6
  PIN b6_c7_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 950.685 32.925 952.140 33.305 ;
        RECT 950.845 30.625 952.140 31.005 ;
        RECT 964.330 30.625 965.640 31.005 ;
        RECT 949.175 29.300 965.185 29.675 ;
        RECT 950.855 25.125 952.160 25.505 ;
        RECT 964.195 25.125 965.660 25.505 ;
        RECT 950.670 23.125 952.160 23.505 ;
      LAYER Metal2 ;
        RECT 950.975 22.415 951.330 33.500 ;
        RECT 964.485 24.845 964.815 31.040 ;
    END
  END b6_c7_not
  PIN b6_c7
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 974.380 33.025 975.660 33.405 ;
        RECT 960.880 30.625 962.065 31.005 ;
        RECT 974.380 30.625 975.395 31.005 ;
        RECT 949.175 27.945 975.405 28.335 ;
        RECT 960.860 25.125 962.220 25.505 ;
        RECT 974.360 25.125 975.540 25.505 ;
        RECT 974.360 23.125 975.435 23.505 ;
      LAYER Metal2 ;
        RECT 961.500 30.990 961.810 31.020 ;
        RECT 961.500 24.890 961.815 30.990 ;
        RECT 975.000 22.895 975.330 33.590 ;
    END
  END b6_c7
  PIN b5_p6
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.615 196.145 1143.745 196.435 ;
        RECT -38.610 73.565 -32.165 73.585 ;
        RECT -38.610 73.300 -5.845 73.565 ;
        RECT -32.500 73.280 -5.845 73.300 ;
        RECT -7.855 72.115 -7.475 72.150 ;
        RECT -29.355 72.010 -28.975 72.050 ;
        RECT -29.425 71.705 -26.590 72.010 ;
        RECT -10.610 71.805 -7.475 72.115 ;
        RECT -7.855 71.770 -7.475 71.805 ;
        RECT -29.355 71.670 -28.975 71.705 ;
        RECT -25.355 63.880 -24.265 64.260 ;
        RECT -12.810 63.880 -11.475 64.260 ;
        RECT -24.870 61.885 -12.020 62.220 ;
        RECT 157.550 53.855 163.995 53.865 ;
        RECT 550.260 53.860 556.705 53.870 ;
        RECT 746.625 53.865 753.070 53.875 ;
        RECT -88.375 53.480 -56.100 53.765 ;
        RECT 157.550 53.580 190.395 53.855 ;
        RECT 163.740 53.570 190.395 53.580 ;
        RECT 353.940 53.815 360.385 53.825 ;
        RECT 353.940 53.540 386.785 53.815 ;
        RECT 550.260 53.585 583.105 53.860 ;
        RECT 746.625 53.590 779.470 53.865 ;
        RECT 556.450 53.575 583.105 53.585 ;
        RECT 752.815 53.580 779.470 53.590 ;
        RECT 943.010 53.850 949.455 53.860 ;
        RECT 1139.335 53.855 1145.780 53.865 ;
        RECT 943.010 53.575 975.855 53.850 ;
        RECT 1139.335 53.580 1172.180 53.855 ;
        RECT 949.200 53.565 975.855 53.575 ;
        RECT 1145.525 53.570 1172.180 53.580 ;
        RECT 360.130 53.530 386.785 53.540 ;
        RECT 188.385 52.405 188.765 52.440 ;
        RECT 581.095 52.410 581.475 52.445 ;
        RECT 777.460 52.415 777.840 52.450 ;
        RECT -58.110 52.315 -57.730 52.350 ;
        RECT -79.610 52.210 -79.230 52.250 ;
        RECT -79.680 51.905 -76.845 52.210 ;
        RECT -60.865 52.005 -57.730 52.315 ;
        RECT 166.885 52.300 167.265 52.340 ;
        RECT -58.110 51.970 -57.730 52.005 ;
        RECT 166.815 51.995 169.650 52.300 ;
        RECT 185.630 52.095 188.765 52.405 ;
        RECT 384.775 52.365 385.155 52.400 ;
        RECT 363.275 52.260 363.655 52.300 ;
        RECT 188.385 52.060 188.765 52.095 ;
        RECT 166.885 51.960 167.265 51.995 ;
        RECT 363.205 51.955 366.040 52.260 ;
        RECT 382.020 52.055 385.155 52.365 ;
        RECT 559.595 52.305 559.975 52.345 ;
        RECT 384.775 52.020 385.155 52.055 ;
        RECT 559.525 52.000 562.360 52.305 ;
        RECT 578.340 52.100 581.475 52.410 ;
        RECT 755.960 52.310 756.340 52.350 ;
        RECT 581.095 52.065 581.475 52.100 ;
        RECT 755.890 52.005 758.725 52.310 ;
        RECT 774.705 52.105 777.840 52.415 ;
        RECT 973.845 52.400 974.225 52.435 ;
        RECT 1170.170 52.405 1170.550 52.440 ;
        RECT 952.345 52.295 952.725 52.335 ;
        RECT 777.460 52.070 777.840 52.105 ;
        RECT 559.595 51.965 559.975 52.000 ;
        RECT 755.960 51.970 756.340 52.005 ;
        RECT 952.275 51.990 955.110 52.295 ;
        RECT 971.090 52.090 974.225 52.400 ;
        RECT 1148.670 52.300 1149.050 52.340 ;
        RECT 973.845 52.055 974.225 52.090 ;
        RECT 1148.600 51.995 1151.435 52.300 ;
        RECT 1167.415 52.095 1170.550 52.405 ;
        RECT 1170.170 52.060 1170.550 52.095 ;
        RECT 952.345 51.955 952.725 51.990 ;
        RECT 1148.670 51.960 1149.050 51.995 ;
        RECT 363.275 51.920 363.655 51.955 ;
        RECT -79.610 51.870 -79.230 51.905 ;
        RECT -75.610 44.080 -74.520 44.460 ;
        RECT -63.065 44.080 -61.730 44.460 ;
        RECT 170.885 44.170 171.975 44.550 ;
        RECT 183.430 44.170 184.765 44.550 ;
        RECT 367.275 44.130 368.365 44.510 ;
        RECT 379.820 44.130 381.155 44.510 ;
        RECT 563.595 44.175 564.685 44.555 ;
        RECT 576.140 44.175 577.475 44.555 ;
        RECT 759.960 44.180 761.050 44.560 ;
        RECT 772.505 44.180 773.840 44.560 ;
        RECT 956.345 44.165 957.435 44.545 ;
        RECT 968.890 44.165 970.225 44.545 ;
        RECT 1152.670 44.170 1153.760 44.550 ;
        RECT 1165.215 44.170 1166.550 44.550 ;
        RECT -75.125 42.085 -62.275 42.420 ;
        RECT 171.370 42.175 184.220 42.510 ;
        RECT 367.760 42.135 380.610 42.470 ;
        RECT 564.080 42.180 576.930 42.515 ;
        RECT 760.445 42.185 773.295 42.520 ;
        RECT 956.830 42.170 969.680 42.505 ;
        RECT 1153.155 42.175 1166.005 42.510 ;
      LAYER Metal2 ;
        RECT -88.080 18.000 -87.790 204.535 ;
        RECT -77.210 51.785 -76.920 53.845 ;
        RECT -74.920 41.870 -74.595 44.635 ;
        RECT -68.340 41.995 -68.050 53.830 ;
        RECT -60.435 51.725 -60.125 54.240 ;
        RECT -62.985 41.870 -62.660 44.635 ;
        RECT -38.340 18.010 -38.000 204.535 ;
        RECT -26.955 71.585 -26.665 73.645 ;
        RECT -24.665 61.670 -24.340 64.435 ;
        RECT -18.085 61.795 -17.795 73.630 ;
        RECT -10.180 71.525 -9.870 74.040 ;
        RECT -12.730 61.670 -12.405 64.435 ;
        RECT 157.830 18.020 158.170 204.545 ;
        RECT 169.285 51.875 169.575 53.935 ;
        RECT 171.575 41.960 171.900 44.725 ;
        RECT 178.155 42.085 178.445 53.920 ;
        RECT 186.060 51.815 186.370 54.330 ;
        RECT 183.510 41.960 183.835 44.725 ;
        RECT 354.220 17.980 354.560 204.505 ;
        RECT 365.675 51.835 365.965 53.895 ;
        RECT 367.965 41.920 368.290 44.685 ;
        RECT 374.545 42.045 374.835 53.880 ;
        RECT 382.450 51.775 382.760 54.290 ;
        RECT 379.900 41.920 380.225 44.685 ;
        RECT 550.540 18.025 550.880 204.550 ;
        RECT 561.995 51.880 562.285 53.940 ;
        RECT 564.285 41.965 564.610 44.730 ;
        RECT 570.865 42.090 571.155 53.925 ;
        RECT 578.770 51.820 579.080 54.335 ;
        RECT 576.220 41.965 576.545 44.730 ;
        RECT 746.905 18.030 747.245 204.555 ;
        RECT 758.360 51.885 758.650 53.945 ;
        RECT 760.650 41.970 760.975 44.735 ;
        RECT 767.230 42.095 767.520 53.930 ;
        RECT 775.135 51.825 775.445 54.340 ;
        RECT 772.585 41.970 772.910 44.735 ;
        RECT 943.290 18.015 943.630 204.540 ;
        RECT 954.745 51.870 955.035 53.930 ;
        RECT 957.035 41.955 957.360 44.720 ;
        RECT 963.615 42.080 963.905 53.915 ;
        RECT 971.520 51.810 971.830 54.325 ;
        RECT 968.970 41.955 969.295 44.720 ;
        RECT 1139.615 18.020 1139.955 204.545 ;
        RECT 1151.070 51.875 1151.360 53.935 ;
        RECT 1153.360 41.960 1153.685 44.725 ;
        RECT 1159.940 42.085 1160.230 53.920 ;
        RECT 1167.845 51.815 1168.155 54.330 ;
        RECT 1165.295 41.960 1165.620 44.725 ;
    END
  END b5_p6
  PIN b5_p7_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.595 194.430 1143.750 194.755 ;
        RECT -21.285 49.985 -20.905 50.030 ;
        RECT -15.785 49.985 -15.405 50.030 ;
        RECT -21.335 49.670 -15.400 49.985 ;
        RECT -21.285 49.650 -20.905 49.670 ;
        RECT -15.785 49.650 -15.405 49.670 ;
        RECT -29.285 42.160 -28.195 42.540 ;
        RECT -7.785 42.495 -7.405 42.540 ;
        RECT -8.520 42.195 -7.210 42.495 ;
        RECT -7.785 42.160 -7.405 42.195 ;
        RECT -32.430 41.645 -5.775 41.650 ;
        RECT -35.155 41.300 -5.775 41.645 ;
        RECT -35.155 41.295 -32.220 41.300 ;
        RECT 174.860 30.265 175.240 30.310 ;
        RECT 180.360 30.265 180.740 30.310 ;
        RECT 567.570 30.270 567.950 30.315 ;
        RECT 573.070 30.270 573.450 30.315 ;
        RECT 763.935 30.275 764.315 30.320 ;
        RECT 769.435 30.275 769.815 30.320 ;
        RECT -71.605 30.095 -71.225 30.140 ;
        RECT -66.105 30.095 -65.725 30.140 ;
        RECT -71.655 29.780 -65.720 30.095 ;
        RECT 174.810 29.950 180.745 30.265 ;
        RECT 371.250 30.225 371.630 30.270 ;
        RECT 376.750 30.225 377.130 30.270 ;
        RECT 174.860 29.930 175.240 29.950 ;
        RECT 180.360 29.930 180.740 29.950 ;
        RECT 371.200 29.910 377.135 30.225 ;
        RECT 567.520 29.955 573.455 30.270 ;
        RECT 763.885 29.960 769.820 30.275 ;
        RECT 960.320 30.260 960.700 30.305 ;
        RECT 965.820 30.260 966.200 30.305 ;
        RECT 1156.645 30.265 1157.025 30.310 ;
        RECT 1162.145 30.265 1162.525 30.310 ;
        RECT 567.570 29.935 567.950 29.955 ;
        RECT 573.070 29.935 573.450 29.955 ;
        RECT 763.935 29.940 764.315 29.960 ;
        RECT 769.435 29.940 769.815 29.960 ;
        RECT 960.270 29.945 966.205 30.260 ;
        RECT 1156.595 29.950 1162.530 30.265 ;
        RECT 960.320 29.925 960.700 29.945 ;
        RECT 965.820 29.925 966.200 29.945 ;
        RECT 1156.645 29.930 1157.025 29.950 ;
        RECT 1162.145 29.930 1162.525 29.950 ;
        RECT 371.250 29.890 371.630 29.910 ;
        RECT 376.750 29.890 377.130 29.910 ;
        RECT -71.605 29.760 -71.225 29.780 ;
        RECT -66.105 29.760 -65.725 29.780 ;
        RECT -79.605 22.270 -78.515 22.650 ;
        RECT -58.105 22.605 -57.725 22.650 ;
        RECT -58.840 22.305 -57.530 22.605 ;
        RECT 166.860 22.440 167.950 22.820 ;
        RECT 188.360 22.775 188.740 22.820 ;
        RECT 187.625 22.475 188.935 22.775 ;
        RECT 188.360 22.440 188.740 22.475 ;
        RECT 363.250 22.400 364.340 22.780 ;
        RECT 384.750 22.735 385.130 22.780 ;
        RECT 384.015 22.435 385.325 22.735 ;
        RECT 559.570 22.445 560.660 22.825 ;
        RECT 581.070 22.780 581.450 22.825 ;
        RECT 580.335 22.480 581.645 22.780 ;
        RECT 581.070 22.445 581.450 22.480 ;
        RECT 755.935 22.450 757.025 22.830 ;
        RECT 777.435 22.785 777.815 22.830 ;
        RECT 776.700 22.485 778.010 22.785 ;
        RECT 777.435 22.450 777.815 22.485 ;
        RECT 952.320 22.435 953.410 22.815 ;
        RECT 973.820 22.770 974.200 22.815 ;
        RECT 973.085 22.470 974.395 22.770 ;
        RECT 973.820 22.435 974.200 22.470 ;
        RECT 1148.645 22.440 1149.735 22.820 ;
        RECT 1170.145 22.775 1170.525 22.820 ;
        RECT 1169.410 22.475 1170.720 22.775 ;
        RECT 1170.145 22.440 1170.525 22.475 ;
        RECT 384.750 22.400 385.130 22.435 ;
        RECT -58.105 22.270 -57.725 22.305 ;
        RECT 752.790 21.935 779.445 21.940 ;
        RECT 556.425 21.930 583.080 21.935 ;
        RECT 163.715 21.925 190.370 21.930 ;
        RECT -82.750 21.755 -56.095 21.760 ;
        RECT -84.915 21.410 -56.095 21.755 ;
        RECT 161.005 21.580 190.370 21.925 ;
        RECT 360.105 21.885 386.760 21.890 ;
        RECT 161.005 21.575 163.940 21.580 ;
        RECT 357.395 21.540 386.760 21.885 ;
        RECT 553.715 21.585 583.080 21.930 ;
        RECT 750.080 21.590 779.445 21.935 ;
        RECT 1145.500 21.925 1172.155 21.930 ;
        RECT 949.175 21.920 975.830 21.925 ;
        RECT 750.080 21.585 753.015 21.590 ;
        RECT 553.715 21.580 556.650 21.585 ;
        RECT 946.465 21.575 975.830 21.920 ;
        RECT 1142.790 21.580 1172.155 21.925 ;
        RECT 1142.790 21.575 1145.725 21.580 ;
        RECT 946.465 21.570 949.400 21.575 ;
        RECT 357.395 21.535 360.330 21.540 ;
        RECT -84.915 21.405 -82.465 21.410 ;
      LAYER Metal2 ;
        RECT -84.740 18.000 -84.380 204.525 ;
        RECT -78.990 21.410 -78.610 22.785 ;
        RECT -69.280 21.120 -68.910 30.220 ;
        RECT -58.735 21.325 -58.400 22.675 ;
        RECT -34.965 17.995 -34.650 204.520 ;
        RECT -28.670 41.300 -28.290 42.675 ;
        RECT -18.960 41.010 -18.590 50.110 ;
        RECT -8.415 41.215 -8.080 42.565 ;
        RECT 161.205 18.005 161.520 204.530 ;
        RECT 167.475 21.580 167.855 22.955 ;
        RECT 177.185 21.290 177.555 30.390 ;
        RECT 187.730 21.495 188.065 22.845 ;
        RECT 357.595 17.965 357.910 204.490 ;
        RECT 363.865 21.540 364.245 22.915 ;
        RECT 373.575 21.250 373.945 30.350 ;
        RECT 384.120 21.455 384.455 22.805 ;
        RECT 553.915 18.010 554.230 204.535 ;
        RECT 560.185 21.585 560.565 22.960 ;
        RECT 569.895 21.295 570.265 30.395 ;
        RECT 580.440 21.500 580.775 22.850 ;
        RECT 750.280 18.015 750.595 204.540 ;
        RECT 756.550 21.590 756.930 22.965 ;
        RECT 766.260 21.300 766.630 30.400 ;
        RECT 776.805 21.505 777.140 22.855 ;
        RECT 946.665 18.000 946.980 204.525 ;
        RECT 952.935 21.575 953.315 22.950 ;
        RECT 962.645 21.285 963.015 30.385 ;
        RECT 973.190 21.490 973.525 22.840 ;
        RECT 1142.990 18.005 1143.305 204.530 ;
        RECT 1149.260 21.580 1149.640 22.955 ;
        RECT 1158.970 21.290 1159.340 30.390 ;
        RECT 1169.515 21.495 1169.850 22.845 ;
    END
  END b5_p7_not
  PIN b5_p7
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.570 195.065 1143.760 195.340 ;
        RECT -32.430 53.840 -5.775 53.845 ;
        RECT -36.440 53.560 -5.775 53.840 ;
        RECT -36.440 53.555 -32.270 53.560 ;
        RECT -7.785 52.395 -7.405 52.430 ;
        RECT -29.285 52.290 -28.905 52.330 ;
        RECT -29.355 51.985 -26.520 52.290 ;
        RECT -10.540 52.085 -7.405 52.395 ;
        RECT -7.785 52.050 -7.405 52.085 ;
        RECT -29.285 51.950 -28.905 51.985 ;
        RECT -25.285 44.160 -24.195 44.540 ;
        RECT -12.740 44.160 -11.405 44.540 ;
        RECT -24.800 42.165 -11.950 42.500 ;
        RECT 752.790 34.130 779.445 34.135 ;
        RECT 556.425 34.125 583.080 34.130 ;
        RECT 163.715 34.120 190.370 34.125 ;
        RECT -82.750 33.950 -56.095 33.955 ;
        RECT -86.195 33.670 -56.095 33.950 ;
        RECT 159.720 33.840 190.370 34.120 ;
        RECT 360.105 34.080 386.760 34.085 ;
        RECT 159.720 33.835 163.890 33.840 ;
        RECT 356.110 33.800 386.760 34.080 ;
        RECT 552.430 33.845 583.080 34.125 ;
        RECT 748.795 33.850 779.445 34.130 ;
        RECT 1145.500 34.120 1172.155 34.125 ;
        RECT 949.175 34.115 975.830 34.120 ;
        RECT 748.795 33.845 752.965 33.850 ;
        RECT 552.430 33.840 556.600 33.845 ;
        RECT 945.180 33.835 975.830 34.115 ;
        RECT 1141.505 33.840 1172.155 34.120 ;
        RECT 1141.505 33.835 1145.675 33.840 ;
        RECT 945.180 33.830 949.350 33.835 ;
        RECT 356.110 33.795 360.280 33.800 ;
        RECT -86.195 33.665 -82.365 33.670 ;
        RECT 188.360 32.675 188.740 32.710 ;
        RECT 581.070 32.680 581.450 32.715 ;
        RECT 777.435 32.685 777.815 32.720 ;
        RECT 166.860 32.570 167.240 32.610 ;
        RECT -58.105 32.505 -57.725 32.540 ;
        RECT -79.605 32.400 -79.225 32.440 ;
        RECT -79.675 32.095 -76.840 32.400 ;
        RECT -60.860 32.195 -57.725 32.505 ;
        RECT 166.790 32.265 169.625 32.570 ;
        RECT 185.605 32.365 188.740 32.675 ;
        RECT 384.750 32.635 385.130 32.670 ;
        RECT 363.250 32.530 363.630 32.570 ;
        RECT 188.360 32.330 188.740 32.365 ;
        RECT 166.860 32.230 167.240 32.265 ;
        RECT 363.180 32.225 366.015 32.530 ;
        RECT 381.995 32.325 385.130 32.635 ;
        RECT 559.570 32.575 559.950 32.615 ;
        RECT 384.750 32.290 385.130 32.325 ;
        RECT 559.500 32.270 562.335 32.575 ;
        RECT 578.315 32.370 581.450 32.680 ;
        RECT 755.935 32.580 756.315 32.620 ;
        RECT 581.070 32.335 581.450 32.370 ;
        RECT 755.865 32.275 758.700 32.580 ;
        RECT 774.680 32.375 777.815 32.685 ;
        RECT 973.820 32.670 974.200 32.705 ;
        RECT 1170.145 32.675 1170.525 32.710 ;
        RECT 952.320 32.565 952.700 32.605 ;
        RECT 777.435 32.340 777.815 32.375 ;
        RECT 559.570 32.235 559.950 32.270 ;
        RECT 755.935 32.240 756.315 32.275 ;
        RECT 952.250 32.260 955.085 32.565 ;
        RECT 971.065 32.360 974.200 32.670 ;
        RECT 1148.645 32.570 1149.025 32.610 ;
        RECT 973.820 32.325 974.200 32.360 ;
        RECT 1148.575 32.265 1151.410 32.570 ;
        RECT 1167.390 32.365 1170.525 32.675 ;
        RECT 1170.145 32.330 1170.525 32.365 ;
        RECT 952.320 32.225 952.700 32.260 ;
        RECT 1148.645 32.230 1149.025 32.265 ;
        RECT -58.105 32.160 -57.725 32.195 ;
        RECT 363.250 32.190 363.630 32.225 ;
        RECT -79.605 32.060 -79.225 32.095 ;
        RECT -75.605 24.270 -74.515 24.650 ;
        RECT -63.060 24.270 -61.725 24.650 ;
        RECT 170.860 24.440 171.950 24.820 ;
        RECT 183.405 24.440 184.740 24.820 ;
        RECT 367.250 24.400 368.340 24.780 ;
        RECT 379.795 24.400 381.130 24.780 ;
        RECT 563.570 24.445 564.660 24.825 ;
        RECT 576.115 24.445 577.450 24.825 ;
        RECT 759.935 24.450 761.025 24.830 ;
        RECT 772.480 24.450 773.815 24.830 ;
        RECT 956.320 24.435 957.410 24.815 ;
        RECT 968.865 24.435 970.200 24.815 ;
        RECT 1152.645 24.440 1153.735 24.820 ;
        RECT 1165.190 24.440 1166.525 24.820 ;
        RECT -75.120 22.275 -62.270 22.610 ;
        RECT 171.345 22.445 184.195 22.780 ;
        RECT 367.735 22.405 380.585 22.740 ;
        RECT 564.055 22.450 576.905 22.785 ;
        RECT 760.420 22.455 773.270 22.790 ;
        RECT 956.805 22.440 969.655 22.775 ;
        RECT 1153.130 22.445 1165.980 22.780 ;
      LAYER Metal2 ;
        RECT -86.025 18.000 -85.575 204.530 ;
        RECT -77.205 31.975 -76.915 34.035 ;
        RECT -74.915 22.060 -74.590 24.825 ;
        RECT -68.335 22.185 -68.045 34.020 ;
        RECT -60.430 31.915 -60.120 34.430 ;
        RECT -62.980 22.060 -62.655 24.825 ;
        RECT -36.210 18.005 -35.890 204.520 ;
        RECT -26.885 51.865 -26.595 53.925 ;
        RECT -24.595 41.950 -24.270 44.715 ;
        RECT -18.015 42.075 -17.725 53.910 ;
        RECT -10.110 51.805 -9.800 54.320 ;
        RECT -12.660 41.950 -12.335 44.715 ;
        RECT 159.960 18.015 160.280 204.530 ;
        RECT 169.260 32.145 169.550 34.205 ;
        RECT 171.550 22.230 171.875 24.995 ;
        RECT 178.130 22.355 178.420 34.190 ;
        RECT 186.035 32.085 186.345 34.600 ;
        RECT 183.485 22.230 183.810 24.995 ;
        RECT 356.350 17.975 356.670 204.490 ;
        RECT 365.650 32.105 365.940 34.165 ;
        RECT 367.940 22.190 368.265 24.955 ;
        RECT 374.520 22.315 374.810 34.150 ;
        RECT 382.425 32.045 382.735 34.560 ;
        RECT 379.875 22.190 380.200 24.955 ;
        RECT 552.670 18.020 552.990 204.535 ;
        RECT 561.970 32.150 562.260 34.210 ;
        RECT 564.260 22.235 564.585 25.000 ;
        RECT 570.840 22.360 571.130 34.195 ;
        RECT 578.745 32.090 579.055 34.605 ;
        RECT 576.195 22.235 576.520 25.000 ;
        RECT 749.035 18.025 749.355 204.540 ;
        RECT 758.335 32.155 758.625 34.215 ;
        RECT 760.625 22.240 760.950 25.005 ;
        RECT 767.205 22.365 767.495 34.200 ;
        RECT 775.110 32.095 775.420 34.610 ;
        RECT 772.560 22.240 772.885 25.005 ;
        RECT 945.420 18.010 945.740 204.525 ;
        RECT 954.720 32.140 955.010 34.200 ;
        RECT 957.010 22.225 957.335 24.990 ;
        RECT 963.590 22.350 963.880 34.185 ;
        RECT 971.495 32.080 971.805 34.595 ;
        RECT 968.945 22.225 969.270 24.990 ;
        RECT 1141.745 18.015 1142.065 204.530 ;
        RECT 1151.045 32.145 1151.335 34.205 ;
        RECT 1153.335 22.230 1153.660 24.995 ;
        RECT 1159.915 22.355 1160.205 34.190 ;
        RECT 1167.820 32.085 1168.130 34.600 ;
        RECT 1165.270 22.230 1165.595 24.995 ;
    END
  END b5_p7
  PIN b5_c7
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 777.995 33.040 779.275 33.420 ;
        RECT 764.495 30.640 765.680 31.020 ;
        RECT 777.995 30.640 779.010 31.020 ;
        RECT 752.790 27.960 779.020 28.350 ;
        RECT 764.475 25.140 765.835 25.520 ;
        RECT 777.975 25.140 779.155 25.520 ;
        RECT 777.975 23.140 779.050 23.520 ;
      LAYER Metal2 ;
        RECT 765.115 31.005 765.425 31.035 ;
        RECT 765.115 24.905 765.430 31.005 ;
        RECT 778.615 22.910 778.945 33.605 ;
    END
  END b5_c7
  PIN b5_c7_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 754.300 32.940 755.755 33.320 ;
        RECT 754.460 30.640 755.755 31.020 ;
        RECT 767.945 30.640 769.255 31.020 ;
        RECT 752.790 29.315 768.800 29.690 ;
        RECT 754.470 25.140 755.775 25.520 ;
        RECT 767.810 25.140 769.275 25.520 ;
        RECT 754.285 23.140 755.775 23.520 ;
      LAYER Metal2 ;
        RECT 754.590 22.430 754.945 33.515 ;
        RECT 768.100 24.860 768.430 31.055 ;
    END
  END b5_c7_not
  PIN b5_c4_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 754.325 92.220 755.780 92.600 ;
        RECT 754.485 89.920 755.780 90.300 ;
        RECT 767.970 89.920 769.280 90.300 ;
        RECT 752.815 88.595 768.825 88.970 ;
        RECT 754.495 84.420 755.800 84.800 ;
        RECT 767.835 84.420 769.300 84.800 ;
        RECT 754.310 82.420 755.800 82.800 ;
      LAYER Metal2 ;
        RECT 754.615 81.710 754.970 92.795 ;
        RECT 768.125 84.140 768.455 90.335 ;
    END
  END b5_c4_not
  PIN x4_b0_f
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 867.460 10.880 867.840 11.260 ;
        RECT 865.860 10.365 867.060 10.655 ;
        RECT 858.125 8.195 867.055 8.495 ;
        RECT 866.650 4.590 867.840 4.875 ;
        RECT 865.870 3.925 866.250 4.305 ;
      LAYER Metal2 ;
        RECT 865.910 3.915 866.210 10.725 ;
        RECT 866.700 4.510 867.010 10.700 ;
        RECT 867.495 4.440 867.795 11.270 ;
    END
  END x4_b0_f
  PIN x4_b0_f_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 861.000 11.100 864.410 11.480 ;
        RECT 872.780 10.430 873.160 10.810 ;
        RECT 858.095 7.660 864.435 7.930 ;
        RECT 864.010 6.400 870.400 6.690 ;
        RECT 860.990 4.485 861.370 4.865 ;
        RECT 869.990 3.760 873.170 4.080 ;
      LAYER Metal2 ;
        RECT 861.035 4.430 861.335 11.470 ;
        RECT 864.060 6.300 864.385 11.460 ;
        RECT 870.070 3.700 870.350 6.735 ;
        RECT 872.820 3.655 873.120 10.810 ;
    END
  END x4_b0_f_not
  PIN x3_b0_f
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 671.120 10.880 671.500 11.260 ;
        RECT 669.520 10.365 670.720 10.655 ;
        RECT 661.785 8.195 670.715 8.495 ;
        RECT 670.310 4.590 671.500 4.875 ;
        RECT 669.530 3.925 669.910 4.305 ;
      LAYER Metal2 ;
        RECT 669.570 3.915 669.870 10.725 ;
        RECT 670.360 4.510 670.670 10.700 ;
        RECT 671.155 4.440 671.455 11.270 ;
    END
  END x3_b0_f
  PIN x3_b0_f_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 664.660 11.100 668.070 11.480 ;
        RECT 676.440 10.430 676.820 10.810 ;
        RECT 661.755 7.660 668.095 7.930 ;
        RECT 667.670 6.400 674.060 6.690 ;
        RECT 664.650 4.485 665.030 4.865 ;
        RECT 673.650 3.760 676.830 4.080 ;
      LAYER Metal2 ;
        RECT 664.695 4.430 664.995 11.470 ;
        RECT 667.720 6.300 668.045 11.460 ;
        RECT 673.730 3.700 674.010 6.735 ;
        RECT 676.480 3.655 676.780 10.810 ;
    END
  END x3_b0_f_not
  PIN p11_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 1308.300 89.915 1308.680 90.295 ;
        RECT 1305.225 89.420 1307.850 89.830 ;
        RECT 1307.410 86.980 1315.110 87.255 ;
        RECT 1307.425 83.555 1308.735 83.875 ;
        RECT 1305.235 83.000 1305.615 83.380 ;
      LAYER Metal2 ;
        RECT 1305.275 82.910 1305.575 89.850 ;
        RECT 1307.485 83.485 1307.765 89.845 ;
        RECT 1308.335 83.485 1308.635 90.305 ;
    END
  END p11_not
  PIN p11
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 1301.400 89.925 1301.780 90.305 ;
        RECT 1298.725 89.500 1300.465 89.790 ;
        RECT 1300.080 84.905 1316.100 85.240 ;
        RECT 1300.050 83.585 1301.830 83.875 ;
        RECT 1298.780 82.970 1299.160 83.350 ;
      LAYER Metal2 ;
        RECT 1298.810 82.910 1299.110 89.840 ;
        RECT 1300.120 83.510 1300.420 89.860 ;
        RECT 1301.435 83.540 1301.730 90.365 ;
    END
  END p11
  PIN p12_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 1308.405 70.200 1308.785 70.580 ;
        RECT 1305.330 69.705 1307.955 70.115 ;
        RECT 1307.515 67.265 1315.215 67.540 ;
        RECT 1307.530 63.840 1308.840 64.160 ;
        RECT 1305.340 63.285 1305.720 63.665 ;
      LAYER Metal2 ;
        RECT 1305.380 63.195 1305.680 70.135 ;
        RECT 1307.590 63.770 1307.870 70.130 ;
        RECT 1308.440 63.770 1308.740 70.590 ;
    END
  END p12_not
  PIN p12
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 1301.505 70.210 1301.885 70.590 ;
        RECT 1298.830 69.785 1300.570 70.075 ;
        RECT 1300.185 65.190 1316.205 65.525 ;
        RECT 1300.155 63.870 1301.935 64.160 ;
        RECT 1298.885 63.255 1299.265 63.635 ;
      LAYER Metal2 ;
        RECT 1298.915 63.195 1299.215 70.125 ;
        RECT 1300.225 63.795 1300.525 70.145 ;
        RECT 1301.540 63.825 1301.835 70.650 ;
    END
  END p12
  PIN p13_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 1308.405 50.230 1308.785 50.610 ;
        RECT 1305.330 49.735 1307.955 50.145 ;
        RECT 1307.515 47.295 1315.215 47.570 ;
        RECT 1307.530 43.870 1308.840 44.190 ;
        RECT 1305.340 43.315 1305.720 43.695 ;
      LAYER Metal2 ;
        RECT 1305.380 43.225 1305.680 50.165 ;
        RECT 1307.590 43.800 1307.870 50.160 ;
        RECT 1308.440 43.800 1308.740 50.620 ;
    END
  END p13_not
  PIN p13
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 1301.505 50.240 1301.885 50.620 ;
        RECT 1298.830 49.815 1300.570 50.105 ;
        RECT 1300.185 45.220 1316.205 45.555 ;
        RECT 1300.155 43.900 1301.935 44.190 ;
        RECT 1298.885 43.285 1299.265 43.665 ;
      LAYER Metal2 ;
        RECT 1298.915 43.225 1299.215 50.155 ;
        RECT 1300.225 43.825 1300.525 50.175 ;
        RECT 1301.540 43.855 1301.835 50.680 ;
    END
  END p13
  PIN p14_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 1308.405 30.565 1308.785 30.945 ;
        RECT 1305.330 30.070 1307.955 30.480 ;
        RECT 1307.515 27.630 1315.215 27.905 ;
        RECT 1307.530 24.205 1308.840 24.525 ;
        RECT 1305.340 23.650 1305.720 24.030 ;
      LAYER Metal2 ;
        RECT 1305.380 23.560 1305.680 30.500 ;
        RECT 1307.590 24.135 1307.870 30.495 ;
        RECT 1308.440 24.135 1308.740 30.955 ;
    END
  END p14_not
  PIN p14
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 1301.505 30.575 1301.885 30.955 ;
        RECT 1298.830 30.150 1300.570 30.440 ;
        RECT 1300.185 25.555 1316.205 25.890 ;
        RECT 1300.155 24.235 1301.935 24.525 ;
        RECT 1298.885 23.620 1299.265 24.000 ;
      LAYER Metal2 ;
        RECT 1298.915 23.560 1299.215 30.490 ;
        RECT 1300.225 24.160 1300.525 30.510 ;
        RECT 1301.540 24.190 1301.835 31.015 ;
    END
  END p14
  PIN b7_c4_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1147.035 92.210 1148.490 92.590 ;
        RECT 1147.195 89.910 1148.490 90.290 ;
        RECT 1160.680 89.910 1161.990 90.290 ;
        RECT 1145.525 88.585 1161.535 88.960 ;
        RECT 1147.205 84.410 1148.510 84.790 ;
        RECT 1160.545 84.410 1162.010 84.790 ;
        RECT 1147.020 82.410 1148.510 82.790 ;
      LAYER Metal2 ;
        RECT 1147.325 81.700 1147.680 92.785 ;
        RECT 1160.835 84.130 1161.165 90.325 ;
    END
  END b7_c4_not
  PIN b7_c4
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1170.730 92.310 1172.010 92.690 ;
        RECT 1157.230 89.910 1158.415 90.290 ;
        RECT 1170.730 89.910 1171.745 90.290 ;
        RECT 1145.525 87.230 1171.755 87.620 ;
        RECT 1157.210 84.410 1158.570 84.790 ;
        RECT 1170.710 84.410 1171.890 84.790 ;
        RECT 1170.710 82.410 1171.785 82.790 ;
      LAYER Metal2 ;
        RECT 1157.850 90.275 1158.160 90.305 ;
        RECT 1157.850 84.175 1158.165 90.275 ;
        RECT 1171.350 82.180 1171.680 92.875 ;
    END
  END b7_c4
  PIN b7_c5_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1146.965 72.380 1148.420 72.760 ;
        RECT 1147.125 70.080 1148.420 70.460 ;
        RECT 1160.610 70.080 1161.920 70.460 ;
        RECT 1145.455 68.755 1161.465 69.130 ;
        RECT 1147.135 64.580 1148.440 64.960 ;
        RECT 1160.475 64.580 1161.940 64.960 ;
        RECT 1146.950 62.580 1148.440 62.960 ;
      LAYER Metal2 ;
        RECT 1147.255 61.870 1147.610 72.955 ;
        RECT 1160.765 64.300 1161.095 70.495 ;
    END
  END b7_c5_not
  PIN b7_c5
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1170.660 72.480 1171.940 72.860 ;
        RECT 1157.160 70.080 1158.345 70.460 ;
        RECT 1170.660 70.080 1171.675 70.460 ;
        RECT 1145.455 67.400 1171.685 67.790 ;
        RECT 1157.140 64.580 1158.500 64.960 ;
        RECT 1170.640 64.580 1171.820 64.960 ;
        RECT 1170.640 62.580 1171.715 62.960 ;
      LAYER Metal2 ;
        RECT 1157.780 70.445 1158.090 70.475 ;
        RECT 1157.780 64.345 1158.095 70.445 ;
        RECT 1171.280 62.350 1171.610 73.045 ;
    END
  END b7_c5
  PIN b7_c6_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1147.035 52.660 1148.490 53.040 ;
        RECT 1147.195 50.360 1148.490 50.740 ;
        RECT 1160.680 50.360 1161.990 50.740 ;
        RECT 1145.525 49.035 1161.535 49.410 ;
        RECT 1147.205 44.860 1148.510 45.240 ;
        RECT 1160.545 44.860 1162.010 45.240 ;
        RECT 1147.020 42.860 1148.510 43.240 ;
      LAYER Metal2 ;
        RECT 1147.325 42.150 1147.680 53.235 ;
        RECT 1160.835 44.580 1161.165 50.775 ;
    END
  END b7_c6_not
  PIN b7_c6
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1170.730 52.760 1172.010 53.140 ;
        RECT 1157.230 50.360 1158.415 50.740 ;
        RECT 1170.730 50.360 1171.745 50.740 ;
        RECT 1145.525 47.680 1171.755 48.070 ;
        RECT 1157.210 44.860 1158.570 45.240 ;
        RECT 1170.710 44.860 1171.890 45.240 ;
        RECT 1170.710 42.860 1171.785 43.240 ;
      LAYER Metal2 ;
        RECT 1157.850 50.725 1158.160 50.755 ;
        RECT 1157.850 44.625 1158.165 50.725 ;
        RECT 1171.350 42.630 1171.680 53.325 ;
    END
  END b7_c6
  PIN b7_c7_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1147.010 32.930 1148.465 33.310 ;
        RECT 1147.170 30.630 1148.465 31.010 ;
        RECT 1160.655 30.630 1161.965 31.010 ;
        RECT 1145.500 29.305 1161.510 29.680 ;
        RECT 1147.180 25.130 1148.485 25.510 ;
        RECT 1160.520 25.130 1161.985 25.510 ;
        RECT 1146.995 23.130 1148.485 23.510 ;
      LAYER Metal2 ;
        RECT 1147.300 22.420 1147.655 33.505 ;
        RECT 1160.810 24.850 1161.140 31.045 ;
    END
  END b7_c7_not
  PIN b7_c7
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1170.705 33.030 1171.985 33.410 ;
        RECT 1157.205 30.630 1158.390 31.010 ;
        RECT 1170.705 30.630 1171.720 31.010 ;
        RECT 1145.500 27.950 1171.730 28.340 ;
        RECT 1157.185 25.130 1158.545 25.510 ;
        RECT 1170.685 25.130 1171.865 25.510 ;
        RECT 1170.685 23.130 1171.760 23.510 ;
      LAYER Metal2 ;
        RECT 1157.825 30.995 1158.135 31.025 ;
        RECT 1157.825 24.895 1158.140 30.995 ;
        RECT 1171.325 22.900 1171.655 33.595 ;
    END
  END b7_c7
  PIN x5_b0_f
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 1063.800 10.880 1064.180 11.260 ;
        RECT 1062.200 10.365 1063.400 10.655 ;
        RECT 1054.465 8.195 1063.395 8.495 ;
        RECT 1062.990 4.590 1064.180 4.875 ;
        RECT 1062.210 3.925 1062.590 4.305 ;
      LAYER Metal2 ;
        RECT 1062.250 3.915 1062.550 10.725 ;
        RECT 1063.040 4.510 1063.350 10.700 ;
        RECT 1063.835 4.440 1064.135 11.270 ;
    END
  END x5_b0_f
  PIN x5_b0_f_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 1057.340 11.100 1060.750 11.480 ;
        RECT 1069.120 10.430 1069.500 10.810 ;
        RECT 1054.435 7.660 1060.775 7.930 ;
        RECT 1060.350 6.400 1066.740 6.690 ;
        RECT 1057.330 4.485 1057.710 4.865 ;
        RECT 1066.330 3.760 1069.510 4.080 ;
      LAYER Metal2 ;
        RECT 1057.375 4.430 1057.675 11.470 ;
        RECT 1060.400 6.300 1060.725 11.460 ;
        RECT 1066.410 3.700 1066.690 6.735 ;
        RECT 1069.160 3.655 1069.460 10.810 ;
    END
  END x5_b0_f_not
  PIN x6_b0_f
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 1260.140 10.880 1260.520 11.260 ;
        RECT 1258.540 10.365 1259.740 10.655 ;
        RECT 1250.805 8.195 1259.735 8.495 ;
        RECT 1259.330 4.590 1260.520 4.875 ;
        RECT 1258.550 3.925 1258.930 4.305 ;
      LAYER Metal2 ;
        RECT 1258.590 3.915 1258.890 10.725 ;
        RECT 1259.380 4.510 1259.690 10.700 ;
        RECT 1260.175 4.440 1260.475 11.270 ;
    END
  END x6_b0_f
  PIN x6_b0_f_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 1253.680 11.100 1257.090 11.480 ;
        RECT 1265.460 10.430 1265.840 10.810 ;
        RECT 1250.775 7.660 1257.115 7.930 ;
        RECT 1256.690 6.400 1263.080 6.690 ;
        RECT 1253.670 4.485 1254.050 4.865 ;
        RECT 1262.670 3.760 1265.850 4.080 ;
      LAYER Metal2 ;
        RECT 1253.715 4.430 1254.015 11.470 ;
        RECT 1256.740 6.300 1257.065 11.460 ;
        RECT 1262.750 3.700 1263.030 6.735 ;
        RECT 1265.500 3.655 1265.800 10.810 ;
    END
  END x6_b0_f_not
  PIN b4_q0
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT 534.785 204.215 536.405 204.540 ;
        RECT 559.660 168.230 560.040 168.610 ;
        RECT 581.160 168.230 581.540 168.610 ;
        RECT 556.515 165.885 575.185 165.895 ;
        RECT 535.600 165.575 583.170 165.885 ;
        RECT 535.600 165.560 556.810 165.575 ;
        RECT 567.660 163.115 568.040 163.120 ;
        RECT 565.180 162.750 568.045 163.115 ;
        RECT 573.160 163.095 573.540 163.120 ;
        RECT 573.145 162.775 575.290 163.095 ;
        RECT 567.660 162.740 568.040 162.750 ;
        RECT 573.160 162.740 573.540 162.775 ;
        RECT 559.575 148.515 559.955 148.895 ;
        RECT 581.075 148.515 581.455 148.895 ;
        RECT 535.620 146.180 556.640 146.190 ;
        RECT 535.620 146.170 575.100 146.180 ;
        RECT 535.620 145.865 583.085 146.170 ;
        RECT 556.430 145.860 583.085 145.865 ;
        RECT 567.575 143.400 567.955 143.405 ;
        RECT 565.095 143.035 567.960 143.400 ;
        RECT 573.075 143.380 573.455 143.405 ;
        RECT 573.060 143.060 575.205 143.380 ;
        RECT 567.575 143.025 567.955 143.035 ;
        RECT 573.075 143.025 573.455 143.060 ;
        RECT 559.635 128.710 560.015 129.090 ;
        RECT 581.135 128.710 581.515 129.090 ;
        RECT 535.570 126.375 556.850 126.380 ;
        RECT 535.570 126.365 575.160 126.375 ;
        RECT 535.570 126.055 583.145 126.365 ;
        RECT 567.635 123.595 568.015 123.600 ;
        RECT 565.155 123.230 568.020 123.595 ;
        RECT 573.135 123.575 573.515 123.600 ;
        RECT 573.120 123.255 575.265 123.575 ;
        RECT 567.635 123.220 568.015 123.230 ;
        RECT 573.135 123.220 573.515 123.255 ;
        RECT 559.565 108.940 559.945 109.320 ;
        RECT 581.065 108.940 581.445 109.320 ;
        RECT 535.575 106.605 556.620 106.620 ;
        RECT 535.575 106.595 575.090 106.605 ;
        RECT 535.575 106.295 583.075 106.595 ;
        RECT 556.420 106.285 583.075 106.295 ;
        RECT 567.565 103.825 567.945 103.830 ;
        RECT 565.085 103.460 567.950 103.825 ;
        RECT 573.065 103.805 573.445 103.830 ;
        RECT 573.050 103.485 575.195 103.805 ;
        RECT 567.565 103.450 567.945 103.460 ;
        RECT 573.065 103.450 573.445 103.485 ;
        RECT 559.595 89.215 559.975 89.595 ;
        RECT 581.095 89.215 581.475 89.595 ;
        RECT 535.560 86.880 556.640 86.885 ;
        RECT 535.560 86.870 575.120 86.880 ;
        RECT 535.560 86.560 583.105 86.870 ;
        RECT 567.595 84.100 567.975 84.105 ;
        RECT 565.115 83.735 567.980 84.100 ;
        RECT 573.095 84.080 573.475 84.105 ;
        RECT 573.080 83.760 575.225 84.080 ;
        RECT 567.595 83.725 567.975 83.735 ;
        RECT 573.095 83.725 573.475 83.760 ;
        RECT 559.525 69.385 559.905 69.765 ;
        RECT 581.025 69.385 581.405 69.765 ;
        RECT 535.545 67.040 575.050 67.050 ;
        RECT 535.545 66.730 583.035 67.040 ;
        RECT 535.545 66.725 556.565 66.730 ;
        RECT 567.525 64.270 567.905 64.275 ;
        RECT 565.045 63.905 567.910 64.270 ;
        RECT 573.025 64.250 573.405 64.275 ;
        RECT 573.010 63.930 575.155 64.250 ;
        RECT 567.525 63.895 567.905 63.905 ;
        RECT 573.025 63.895 573.405 63.930 ;
        RECT 559.595 49.665 559.975 50.045 ;
        RECT 581.095 49.665 581.475 50.045 ;
        RECT 535.655 47.330 556.705 47.340 ;
        RECT 535.655 47.320 575.120 47.330 ;
        RECT 535.655 47.015 583.105 47.320 ;
        RECT 556.450 47.010 583.105 47.015 ;
        RECT 567.595 44.550 567.975 44.555 ;
        RECT 565.115 44.185 567.980 44.550 ;
        RECT 573.095 44.530 573.475 44.555 ;
        RECT 573.080 44.210 575.225 44.530 ;
        RECT 567.595 44.175 567.975 44.185 ;
        RECT 573.095 44.175 573.475 44.210 ;
        RECT 559.570 29.935 559.950 30.315 ;
        RECT 581.070 29.935 581.450 30.315 ;
        RECT 556.425 27.595 575.095 27.600 ;
        RECT 535.590 27.590 575.095 27.595 ;
        RECT 535.590 27.280 583.080 27.590 ;
        RECT 535.590 27.270 556.570 27.280 ;
        RECT 567.570 24.820 567.950 24.825 ;
        RECT 565.090 24.455 567.955 24.820 ;
        RECT 573.070 24.800 573.450 24.825 ;
        RECT 573.055 24.480 575.200 24.800 ;
        RECT 567.570 24.445 567.950 24.455 ;
        RECT 573.070 24.445 573.450 24.480 ;
      LAYER Metal2 ;
        RECT 535.810 17.845 536.205 204.540 ;
        RECT 559.610 165.575 560.060 168.565 ;
        RECT 565.335 162.565 565.740 165.895 ;
        RECT 574.770 162.620 575.220 165.895 ;
        RECT 581.125 165.575 581.575 168.585 ;
        RECT 559.525 145.860 559.975 148.850 ;
        RECT 565.250 142.850 565.655 146.180 ;
        RECT 574.685 142.905 575.135 146.180 ;
        RECT 581.040 145.860 581.490 148.870 ;
        RECT 559.585 126.055 560.035 129.045 ;
        RECT 565.310 123.045 565.715 126.375 ;
        RECT 574.745 123.100 575.195 126.375 ;
        RECT 581.100 126.055 581.550 129.065 ;
        RECT 559.515 106.285 559.965 109.275 ;
        RECT 565.240 103.275 565.645 106.605 ;
        RECT 574.675 103.330 575.125 106.605 ;
        RECT 581.030 106.285 581.480 109.295 ;
        RECT 559.545 86.560 559.995 89.550 ;
        RECT 565.270 83.550 565.675 86.880 ;
        RECT 574.705 83.605 575.155 86.880 ;
        RECT 581.060 86.560 581.510 89.570 ;
        RECT 559.475 66.730 559.925 69.720 ;
        RECT 565.200 63.720 565.605 67.050 ;
        RECT 574.635 63.775 575.085 67.050 ;
        RECT 580.990 66.730 581.440 69.740 ;
        RECT 559.545 47.010 559.995 50.000 ;
        RECT 565.270 44.000 565.675 47.330 ;
        RECT 574.705 44.055 575.155 47.330 ;
        RECT 581.060 47.010 581.510 50.020 ;
        RECT 559.520 27.280 559.970 30.270 ;
        RECT 565.245 24.270 565.650 27.600 ;
        RECT 574.680 24.325 575.130 27.600 ;
        RECT 581.035 27.280 581.485 30.290 ;
    END
  END b4_q0
  PIN b4_q0_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT 534.770 203.640 537.330 203.945 ;
        RECT 563.660 168.230 564.040 168.610 ;
        RECT 577.160 168.230 577.540 168.610 ;
        RECT 556.515 164.895 583.170 164.905 ;
        RECT 536.760 164.635 583.170 164.895 ;
        RECT 536.760 164.625 556.755 164.635 ;
        RECT 559.660 163.085 560.040 163.120 ;
        RECT 581.160 163.100 581.540 163.120 ;
        RECT 559.395 162.775 562.405 163.085 ;
        RECT 578.695 162.780 581.605 163.100 ;
        RECT 559.660 162.740 560.040 162.775 ;
        RECT 581.160 162.740 581.540 162.780 ;
        RECT 563.575 148.515 563.955 148.895 ;
        RECT 577.075 148.515 577.455 148.895 ;
        RECT 536.780 145.190 556.585 145.200 ;
        RECT 536.780 144.930 583.085 145.190 ;
        RECT 556.430 144.920 583.085 144.930 ;
        RECT 559.575 143.370 559.955 143.405 ;
        RECT 581.075 143.385 581.455 143.405 ;
        RECT 559.310 143.060 562.320 143.370 ;
        RECT 578.610 143.065 581.520 143.385 ;
        RECT 559.575 143.025 559.955 143.060 ;
        RECT 581.075 143.025 581.455 143.065 ;
        RECT 563.635 128.710 564.015 129.090 ;
        RECT 577.135 128.710 577.515 129.090 ;
        RECT 536.730 125.385 556.815 125.390 ;
        RECT 536.730 125.120 583.145 125.385 ;
        RECT 556.490 125.115 583.145 125.120 ;
        RECT 559.635 123.565 560.015 123.600 ;
        RECT 581.135 123.580 581.515 123.600 ;
        RECT 559.370 123.255 562.380 123.565 ;
        RECT 578.670 123.260 581.580 123.580 ;
        RECT 559.635 123.220 560.015 123.255 ;
        RECT 581.135 123.220 581.515 123.260 ;
        RECT 563.565 108.940 563.945 109.320 ;
        RECT 577.065 108.940 577.445 109.320 ;
        RECT 536.735 105.615 556.640 105.630 ;
        RECT 536.735 105.360 583.075 105.615 ;
        RECT 556.420 105.345 583.075 105.360 ;
        RECT 559.565 103.795 559.945 103.830 ;
        RECT 581.065 103.810 581.445 103.830 ;
        RECT 559.300 103.485 562.310 103.795 ;
        RECT 578.600 103.490 581.510 103.810 ;
        RECT 559.565 103.450 559.945 103.485 ;
        RECT 581.065 103.450 581.445 103.490 ;
        RECT 563.595 89.215 563.975 89.595 ;
        RECT 577.095 89.215 577.475 89.595 ;
        RECT 536.720 85.890 556.695 85.895 ;
        RECT 536.720 85.625 583.105 85.890 ;
        RECT 556.450 85.620 583.105 85.625 ;
        RECT 559.595 84.070 559.975 84.105 ;
        RECT 581.095 84.085 581.475 84.105 ;
        RECT 559.330 83.760 562.340 84.070 ;
        RECT 578.630 83.765 581.540 84.085 ;
        RECT 559.595 83.725 559.975 83.760 ;
        RECT 581.095 83.725 581.475 83.765 ;
        RECT 563.525 69.385 563.905 69.765 ;
        RECT 577.025 69.385 577.405 69.765 ;
        RECT 536.700 65.790 583.035 66.060 ;
        RECT 559.525 64.240 559.905 64.275 ;
        RECT 581.025 64.255 581.405 64.275 ;
        RECT 559.260 63.930 562.270 64.240 ;
        RECT 578.560 63.935 581.470 64.255 ;
        RECT 559.525 63.895 559.905 63.930 ;
        RECT 581.025 63.895 581.405 63.935 ;
        RECT 563.595 49.665 563.975 50.045 ;
        RECT 577.095 49.665 577.475 50.045 ;
        RECT 536.815 46.340 556.705 46.350 ;
        RECT 536.815 46.080 583.105 46.340 ;
        RECT 556.450 46.070 583.105 46.080 ;
        RECT 559.595 44.520 559.975 44.555 ;
        RECT 581.095 44.535 581.475 44.555 ;
        RECT 559.330 44.210 562.340 44.520 ;
        RECT 578.630 44.215 581.540 44.535 ;
        RECT 559.595 44.175 559.975 44.210 ;
        RECT 581.095 44.175 581.475 44.215 ;
        RECT 563.570 29.935 563.950 30.315 ;
        RECT 577.070 29.935 577.450 30.315 ;
        RECT 556.425 26.605 583.080 26.610 ;
        RECT 536.750 26.340 583.080 26.605 ;
        RECT 536.750 26.335 556.650 26.340 ;
        RECT 559.570 24.790 559.950 24.825 ;
        RECT 581.070 24.805 581.450 24.825 ;
        RECT 559.305 24.480 562.315 24.790 ;
        RECT 578.605 24.485 581.515 24.805 ;
        RECT 559.570 24.445 559.950 24.480 ;
        RECT 581.070 24.445 581.450 24.485 ;
      LAYER Metal2 ;
        RECT 536.915 17.930 537.255 204.530 ;
        RECT 562.010 162.590 562.305 164.960 ;
        RECT 563.620 164.635 564.070 168.600 ;
        RECT 577.150 164.635 577.550 168.575 ;
        RECT 578.800 162.625 579.215 165.015 ;
        RECT 561.925 142.875 562.220 145.245 ;
        RECT 563.535 144.920 563.985 148.885 ;
        RECT 577.065 144.920 577.465 148.860 ;
        RECT 578.715 142.910 579.130 145.300 ;
        RECT 561.985 123.070 562.280 125.440 ;
        RECT 563.595 125.115 564.045 129.080 ;
        RECT 577.125 125.115 577.525 129.055 ;
        RECT 578.775 123.105 579.190 125.495 ;
        RECT 561.915 103.300 562.210 105.670 ;
        RECT 563.525 105.345 563.975 109.310 ;
        RECT 577.055 105.345 577.455 109.285 ;
        RECT 578.705 103.335 579.120 105.725 ;
        RECT 561.945 83.575 562.240 85.945 ;
        RECT 563.555 85.620 564.005 89.585 ;
        RECT 577.085 85.620 577.485 89.560 ;
        RECT 578.735 83.610 579.150 86.000 ;
        RECT 561.875 63.745 562.170 66.115 ;
        RECT 563.485 65.790 563.935 69.755 ;
        RECT 577.015 65.790 577.415 69.730 ;
        RECT 578.665 63.780 579.080 66.170 ;
        RECT 561.945 44.025 562.240 46.395 ;
        RECT 563.555 46.070 564.005 50.035 ;
        RECT 577.085 46.070 577.485 50.010 ;
        RECT 578.735 44.060 579.150 46.450 ;
        RECT 561.920 24.295 562.215 26.665 ;
        RECT 563.530 26.340 563.980 30.305 ;
        RECT 577.060 26.340 577.460 30.280 ;
        RECT 578.710 24.330 579.125 26.720 ;
    END
  END b4_q0_not
  PIN b3_q0
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT 338.465 204.170 340.085 204.495 ;
        RECT 363.340 168.185 363.720 168.565 ;
        RECT 384.840 168.185 385.220 168.565 ;
        RECT 360.195 165.840 378.865 165.850 ;
        RECT 339.280 165.530 386.850 165.840 ;
        RECT 339.280 165.515 360.490 165.530 ;
        RECT 371.340 163.070 371.720 163.075 ;
        RECT 368.860 162.705 371.725 163.070 ;
        RECT 376.840 163.050 377.220 163.075 ;
        RECT 376.825 162.730 378.970 163.050 ;
        RECT 371.340 162.695 371.720 162.705 ;
        RECT 376.840 162.695 377.220 162.730 ;
        RECT 363.255 148.470 363.635 148.850 ;
        RECT 384.755 148.470 385.135 148.850 ;
        RECT 339.300 146.135 360.320 146.145 ;
        RECT 339.300 146.125 378.780 146.135 ;
        RECT 339.300 145.820 386.765 146.125 ;
        RECT 360.110 145.815 386.765 145.820 ;
        RECT 371.255 143.355 371.635 143.360 ;
        RECT 368.775 142.990 371.640 143.355 ;
        RECT 376.755 143.335 377.135 143.360 ;
        RECT 376.740 143.015 378.885 143.335 ;
        RECT 371.255 142.980 371.635 142.990 ;
        RECT 376.755 142.980 377.135 143.015 ;
        RECT 363.315 128.665 363.695 129.045 ;
        RECT 384.815 128.665 385.195 129.045 ;
        RECT 339.250 126.330 360.530 126.335 ;
        RECT 339.250 126.320 378.840 126.330 ;
        RECT 339.250 126.010 386.825 126.320 ;
        RECT 371.315 123.550 371.695 123.555 ;
        RECT 368.835 123.185 371.700 123.550 ;
        RECT 376.815 123.530 377.195 123.555 ;
        RECT 376.800 123.210 378.945 123.530 ;
        RECT 371.315 123.175 371.695 123.185 ;
        RECT 376.815 123.175 377.195 123.210 ;
        RECT 363.245 108.895 363.625 109.275 ;
        RECT 384.745 108.895 385.125 109.275 ;
        RECT 339.255 106.560 360.300 106.575 ;
        RECT 339.255 106.550 378.770 106.560 ;
        RECT 339.255 106.250 386.755 106.550 ;
        RECT 360.100 106.240 386.755 106.250 ;
        RECT 371.245 103.780 371.625 103.785 ;
        RECT 368.765 103.415 371.630 103.780 ;
        RECT 376.745 103.760 377.125 103.785 ;
        RECT 376.730 103.440 378.875 103.760 ;
        RECT 371.245 103.405 371.625 103.415 ;
        RECT 376.745 103.405 377.125 103.440 ;
        RECT 363.275 89.170 363.655 89.550 ;
        RECT 384.775 89.170 385.155 89.550 ;
        RECT 339.240 86.835 360.320 86.840 ;
        RECT 339.240 86.825 378.800 86.835 ;
        RECT 339.240 86.515 386.785 86.825 ;
        RECT 371.275 84.055 371.655 84.060 ;
        RECT 368.795 83.690 371.660 84.055 ;
        RECT 376.775 84.035 377.155 84.060 ;
        RECT 376.760 83.715 378.905 84.035 ;
        RECT 371.275 83.680 371.655 83.690 ;
        RECT 376.775 83.680 377.155 83.715 ;
        RECT 363.205 69.340 363.585 69.720 ;
        RECT 384.705 69.340 385.085 69.720 ;
        RECT 339.225 66.995 378.730 67.005 ;
        RECT 339.225 66.685 386.715 66.995 ;
        RECT 339.225 66.680 360.245 66.685 ;
        RECT 371.205 64.225 371.585 64.230 ;
        RECT 368.725 63.860 371.590 64.225 ;
        RECT 376.705 64.205 377.085 64.230 ;
        RECT 376.690 63.885 378.835 64.205 ;
        RECT 371.205 63.850 371.585 63.860 ;
        RECT 376.705 63.850 377.085 63.885 ;
        RECT 363.275 49.620 363.655 50.000 ;
        RECT 384.775 49.620 385.155 50.000 ;
        RECT 339.335 47.285 360.385 47.295 ;
        RECT 339.335 47.275 378.800 47.285 ;
        RECT 339.335 46.970 386.785 47.275 ;
        RECT 360.130 46.965 386.785 46.970 ;
        RECT 371.275 44.505 371.655 44.510 ;
        RECT 368.795 44.140 371.660 44.505 ;
        RECT 376.775 44.485 377.155 44.510 ;
        RECT 376.760 44.165 378.905 44.485 ;
        RECT 371.275 44.130 371.655 44.140 ;
        RECT 376.775 44.130 377.155 44.165 ;
        RECT 363.250 29.890 363.630 30.270 ;
        RECT 384.750 29.890 385.130 30.270 ;
        RECT 360.105 27.550 378.775 27.555 ;
        RECT 339.270 27.545 378.775 27.550 ;
        RECT 339.270 27.235 386.760 27.545 ;
        RECT 339.270 27.225 360.250 27.235 ;
        RECT 371.250 24.775 371.630 24.780 ;
        RECT 368.770 24.410 371.635 24.775 ;
        RECT 376.750 24.755 377.130 24.780 ;
        RECT 376.735 24.435 378.880 24.755 ;
        RECT 371.250 24.400 371.630 24.410 ;
        RECT 376.750 24.400 377.130 24.435 ;
      LAYER Metal2 ;
        RECT 339.490 17.800 339.885 204.495 ;
        RECT 363.290 165.530 363.740 168.520 ;
        RECT 369.015 162.520 369.420 165.850 ;
        RECT 378.450 162.575 378.900 165.850 ;
        RECT 384.805 165.530 385.255 168.540 ;
        RECT 363.205 145.815 363.655 148.805 ;
        RECT 368.930 142.805 369.335 146.135 ;
        RECT 378.365 142.860 378.815 146.135 ;
        RECT 384.720 145.815 385.170 148.825 ;
        RECT 363.265 126.010 363.715 129.000 ;
        RECT 368.990 123.000 369.395 126.330 ;
        RECT 378.425 123.055 378.875 126.330 ;
        RECT 384.780 126.010 385.230 129.020 ;
        RECT 363.195 106.240 363.645 109.230 ;
        RECT 368.920 103.230 369.325 106.560 ;
        RECT 378.355 103.285 378.805 106.560 ;
        RECT 384.710 106.240 385.160 109.250 ;
        RECT 363.225 86.515 363.675 89.505 ;
        RECT 368.950 83.505 369.355 86.835 ;
        RECT 378.385 83.560 378.835 86.835 ;
        RECT 384.740 86.515 385.190 89.525 ;
        RECT 363.155 66.685 363.605 69.675 ;
        RECT 368.880 63.675 369.285 67.005 ;
        RECT 378.315 63.730 378.765 67.005 ;
        RECT 384.670 66.685 385.120 69.695 ;
        RECT 363.225 46.965 363.675 49.955 ;
        RECT 368.950 43.955 369.355 47.285 ;
        RECT 378.385 44.010 378.835 47.285 ;
        RECT 384.740 46.965 385.190 49.975 ;
        RECT 363.200 27.235 363.650 30.225 ;
        RECT 368.925 24.225 369.330 27.555 ;
        RECT 378.360 24.280 378.810 27.555 ;
        RECT 384.715 27.235 385.165 30.245 ;
    END
  END b3_q0
  PIN b3_q0_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT 338.450 203.595 341.010 203.900 ;
        RECT 367.340 168.185 367.720 168.565 ;
        RECT 380.840 168.185 381.220 168.565 ;
        RECT 360.195 164.850 386.850 164.860 ;
        RECT 340.440 164.590 386.850 164.850 ;
        RECT 340.440 164.580 360.435 164.590 ;
        RECT 363.340 163.040 363.720 163.075 ;
        RECT 384.840 163.055 385.220 163.075 ;
        RECT 363.075 162.730 366.085 163.040 ;
        RECT 382.375 162.735 385.285 163.055 ;
        RECT 363.340 162.695 363.720 162.730 ;
        RECT 384.840 162.695 385.220 162.735 ;
        RECT 367.255 148.470 367.635 148.850 ;
        RECT 380.755 148.470 381.135 148.850 ;
        RECT 340.460 145.145 360.265 145.155 ;
        RECT 340.460 144.885 386.765 145.145 ;
        RECT 360.110 144.875 386.765 144.885 ;
        RECT 363.255 143.325 363.635 143.360 ;
        RECT 384.755 143.340 385.135 143.360 ;
        RECT 362.990 143.015 366.000 143.325 ;
        RECT 382.290 143.020 385.200 143.340 ;
        RECT 363.255 142.980 363.635 143.015 ;
        RECT 384.755 142.980 385.135 143.020 ;
        RECT 367.315 128.665 367.695 129.045 ;
        RECT 380.815 128.665 381.195 129.045 ;
        RECT 340.410 125.340 360.495 125.345 ;
        RECT 340.410 125.075 386.825 125.340 ;
        RECT 360.170 125.070 386.825 125.075 ;
        RECT 363.315 123.520 363.695 123.555 ;
        RECT 384.815 123.535 385.195 123.555 ;
        RECT 363.050 123.210 366.060 123.520 ;
        RECT 382.350 123.215 385.260 123.535 ;
        RECT 363.315 123.175 363.695 123.210 ;
        RECT 384.815 123.175 385.195 123.215 ;
        RECT 367.245 108.895 367.625 109.275 ;
        RECT 380.745 108.895 381.125 109.275 ;
        RECT 340.415 105.570 360.320 105.585 ;
        RECT 340.415 105.315 386.755 105.570 ;
        RECT 360.100 105.300 386.755 105.315 ;
        RECT 363.245 103.750 363.625 103.785 ;
        RECT 384.745 103.765 385.125 103.785 ;
        RECT 362.980 103.440 365.990 103.750 ;
        RECT 382.280 103.445 385.190 103.765 ;
        RECT 363.245 103.405 363.625 103.440 ;
        RECT 384.745 103.405 385.125 103.445 ;
        RECT 367.275 89.170 367.655 89.550 ;
        RECT 380.775 89.170 381.155 89.550 ;
        RECT 340.400 85.845 360.375 85.850 ;
        RECT 340.400 85.580 386.785 85.845 ;
        RECT 360.130 85.575 386.785 85.580 ;
        RECT 363.275 84.025 363.655 84.060 ;
        RECT 384.775 84.040 385.155 84.060 ;
        RECT 363.010 83.715 366.020 84.025 ;
        RECT 382.310 83.720 385.220 84.040 ;
        RECT 363.275 83.680 363.655 83.715 ;
        RECT 384.775 83.680 385.155 83.720 ;
        RECT 367.205 69.340 367.585 69.720 ;
        RECT 380.705 69.340 381.085 69.720 ;
        RECT 340.380 65.745 386.715 66.015 ;
        RECT 363.205 64.195 363.585 64.230 ;
        RECT 384.705 64.210 385.085 64.230 ;
        RECT 362.940 63.885 365.950 64.195 ;
        RECT 382.240 63.890 385.150 64.210 ;
        RECT 363.205 63.850 363.585 63.885 ;
        RECT 384.705 63.850 385.085 63.890 ;
        RECT 367.275 49.620 367.655 50.000 ;
        RECT 380.775 49.620 381.155 50.000 ;
        RECT 340.495 46.295 360.385 46.305 ;
        RECT 340.495 46.035 386.785 46.295 ;
        RECT 360.130 46.025 386.785 46.035 ;
        RECT 363.275 44.475 363.655 44.510 ;
        RECT 384.775 44.490 385.155 44.510 ;
        RECT 363.010 44.165 366.020 44.475 ;
        RECT 382.310 44.170 385.220 44.490 ;
        RECT 363.275 44.130 363.655 44.165 ;
        RECT 384.775 44.130 385.155 44.170 ;
        RECT 367.250 29.890 367.630 30.270 ;
        RECT 380.750 29.890 381.130 30.270 ;
        RECT 360.105 26.560 386.760 26.565 ;
        RECT 340.430 26.295 386.760 26.560 ;
        RECT 340.430 26.290 360.330 26.295 ;
        RECT 363.250 24.745 363.630 24.780 ;
        RECT 384.750 24.760 385.130 24.780 ;
        RECT 362.985 24.435 365.995 24.745 ;
        RECT 382.285 24.440 385.195 24.760 ;
        RECT 363.250 24.400 363.630 24.435 ;
        RECT 384.750 24.400 385.130 24.440 ;
      LAYER Metal2 ;
        RECT 340.595 17.885 340.935 204.485 ;
        RECT 365.690 162.545 365.985 164.915 ;
        RECT 367.300 164.590 367.750 168.555 ;
        RECT 380.830 164.590 381.230 168.530 ;
        RECT 382.480 162.580 382.895 164.970 ;
        RECT 365.605 142.830 365.900 145.200 ;
        RECT 367.215 144.875 367.665 148.840 ;
        RECT 380.745 144.875 381.145 148.815 ;
        RECT 382.395 142.865 382.810 145.255 ;
        RECT 365.665 123.025 365.960 125.395 ;
        RECT 367.275 125.070 367.725 129.035 ;
        RECT 380.805 125.070 381.205 129.010 ;
        RECT 382.455 123.060 382.870 125.450 ;
        RECT 365.595 103.255 365.890 105.625 ;
        RECT 367.205 105.300 367.655 109.265 ;
        RECT 380.735 105.300 381.135 109.240 ;
        RECT 382.385 103.290 382.800 105.680 ;
        RECT 365.625 83.530 365.920 85.900 ;
        RECT 367.235 85.575 367.685 89.540 ;
        RECT 380.765 85.575 381.165 89.515 ;
        RECT 382.415 83.565 382.830 85.955 ;
        RECT 365.555 63.700 365.850 66.070 ;
        RECT 367.165 65.745 367.615 69.710 ;
        RECT 380.695 65.745 381.095 69.685 ;
        RECT 382.345 63.735 382.760 66.125 ;
        RECT 365.625 43.980 365.920 46.350 ;
        RECT 367.235 46.025 367.685 49.990 ;
        RECT 380.765 46.025 381.165 49.965 ;
        RECT 382.415 44.015 382.830 46.405 ;
        RECT 365.600 24.250 365.895 26.620 ;
        RECT 367.210 26.295 367.660 30.260 ;
        RECT 380.740 26.295 381.140 30.235 ;
        RECT 382.390 24.285 382.805 26.675 ;
    END
  END b3_q0_not
  PIN p2_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 326.630 168.850 327.010 169.230 ;
        RECT 323.555 168.355 326.180 168.765 ;
        RECT 325.740 165.915 333.440 166.190 ;
        RECT 325.755 162.490 327.065 162.810 ;
        RECT 323.565 161.935 323.945 162.315 ;
      LAYER Metal2 ;
        RECT 323.605 161.845 323.905 168.785 ;
        RECT 325.815 162.420 326.095 168.780 ;
        RECT 326.665 162.420 326.965 169.240 ;
    END
  END p2_not
  PIN p2
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 319.730 168.860 320.110 169.240 ;
        RECT 317.055 168.435 318.795 168.725 ;
        RECT 318.410 163.840 334.430 164.175 ;
        RECT 318.380 162.520 320.160 162.810 ;
        RECT 317.110 161.905 317.490 162.285 ;
      LAYER Metal2 ;
        RECT 317.140 161.845 317.440 168.775 ;
        RECT 318.450 162.445 318.750 168.795 ;
        RECT 319.765 162.475 320.060 169.300 ;
    END
  END p2
  PIN p3_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 523.030 168.800 523.410 169.180 ;
        RECT 519.955 168.305 522.580 168.715 ;
        RECT 522.140 165.865 529.840 166.140 ;
        RECT 522.155 162.440 523.465 162.760 ;
        RECT 519.965 161.885 520.345 162.265 ;
      LAYER Metal2 ;
        RECT 520.005 161.795 520.305 168.735 ;
        RECT 522.215 162.370 522.495 168.730 ;
        RECT 523.065 162.370 523.365 169.190 ;
    END
  END p3_not
  PIN p3
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 516.130 168.810 516.510 169.190 ;
        RECT 513.455 168.385 515.195 168.675 ;
        RECT 514.810 163.790 530.830 164.125 ;
        RECT 514.780 162.470 516.560 162.760 ;
        RECT 513.510 161.855 513.890 162.235 ;
      LAYER Metal2 ;
        RECT 513.540 161.795 513.840 168.725 ;
        RECT 514.850 162.395 515.150 168.745 ;
        RECT 516.165 162.425 516.460 169.250 ;
    END
  END p3
  PIN b3_c0_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 361.705 171.185 363.160 171.565 ;
        RECT 361.865 168.885 363.160 169.265 ;
        RECT 375.350 168.885 376.660 169.265 ;
        RECT 360.195 167.560 376.205 167.935 ;
        RECT 361.875 163.385 363.180 163.765 ;
        RECT 375.215 163.385 376.680 163.765 ;
        RECT 361.690 161.385 363.180 161.765 ;
      LAYER Metal2 ;
        RECT 361.995 160.675 362.350 171.760 ;
        RECT 375.505 163.105 375.835 169.300 ;
    END
  END b3_c0_not
  PIN b3_c1_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 361.620 151.470 363.075 151.850 ;
        RECT 361.780 149.170 363.075 149.550 ;
        RECT 375.265 149.170 376.575 149.550 ;
        RECT 360.110 147.845 376.120 148.220 ;
        RECT 361.790 143.670 363.095 144.050 ;
        RECT 375.130 143.670 376.595 144.050 ;
        RECT 361.605 141.670 363.095 142.050 ;
      LAYER Metal2 ;
        RECT 361.910 140.960 362.265 152.045 ;
        RECT 375.420 143.390 375.750 149.585 ;
    END
  END b3_c1_not
  PIN b3_c0
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 385.400 171.285 386.680 171.665 ;
        RECT 371.900 168.885 373.085 169.265 ;
        RECT 385.400 168.885 386.415 169.265 ;
        RECT 360.195 166.205 386.425 166.595 ;
        RECT 371.880 163.385 373.240 163.765 ;
        RECT 385.380 163.385 386.560 163.765 ;
        RECT 385.380 161.385 386.455 161.765 ;
      LAYER Metal2 ;
        RECT 372.520 169.250 372.830 169.280 ;
        RECT 372.520 163.150 372.835 169.250 ;
        RECT 386.020 161.155 386.350 171.850 ;
    END
  END b3_c0
  PIN b3_c1
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 385.315 151.570 386.595 151.950 ;
        RECT 371.815 149.170 373.000 149.550 ;
        RECT 385.315 149.170 386.330 149.550 ;
        RECT 360.110 146.490 386.340 146.880 ;
        RECT 371.795 143.670 373.155 144.050 ;
        RECT 385.295 143.670 386.475 144.050 ;
        RECT 385.295 141.670 386.370 142.050 ;
      LAYER Metal2 ;
        RECT 372.435 149.535 372.745 149.565 ;
        RECT 372.435 143.435 372.750 149.535 ;
        RECT 385.935 141.440 386.265 152.135 ;
    END
  END b3_c1
  PIN b3_c2_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 361.680 131.665 363.135 132.045 ;
        RECT 361.840 129.365 363.135 129.745 ;
        RECT 375.325 129.365 376.635 129.745 ;
        RECT 360.170 128.040 376.180 128.415 ;
        RECT 361.850 123.865 363.155 124.245 ;
        RECT 375.190 123.865 376.655 124.245 ;
        RECT 361.665 121.865 363.155 122.245 ;
      LAYER Metal2 ;
        RECT 361.970 121.155 362.325 132.240 ;
        RECT 375.480 123.585 375.810 129.780 ;
    END
  END b3_c2_not
  PIN b3_c2
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 385.375 131.765 386.655 132.145 ;
        RECT 371.875 129.365 373.060 129.745 ;
        RECT 385.375 129.365 386.390 129.745 ;
        RECT 360.170 126.685 386.400 127.075 ;
        RECT 371.855 123.865 373.215 124.245 ;
        RECT 385.355 123.865 386.535 124.245 ;
        RECT 385.355 121.865 386.430 122.245 ;
      LAYER Metal2 ;
        RECT 372.495 129.730 372.805 129.760 ;
        RECT 372.495 123.630 372.810 129.730 ;
        RECT 385.995 121.635 386.325 132.330 ;
    END
  END b3_c2
  PIN b3_c3_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 361.610 111.895 363.065 112.275 ;
        RECT 361.770 109.595 363.065 109.975 ;
        RECT 375.255 109.595 376.565 109.975 ;
        RECT 360.100 108.270 376.110 108.645 ;
        RECT 361.780 104.095 363.085 104.475 ;
        RECT 375.120 104.095 376.585 104.475 ;
        RECT 361.595 102.095 363.085 102.475 ;
      LAYER Metal2 ;
        RECT 361.900 101.385 362.255 112.470 ;
        RECT 375.410 103.815 375.740 110.010 ;
    END
  END b3_c3_not
  PIN b3_c3
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 385.305 111.995 386.585 112.375 ;
        RECT 371.805 109.595 372.990 109.975 ;
        RECT 385.305 109.595 386.320 109.975 ;
        RECT 360.100 106.915 386.330 107.305 ;
        RECT 371.785 104.095 373.145 104.475 ;
        RECT 385.285 104.095 386.465 104.475 ;
        RECT 385.285 102.095 386.360 102.475 ;
      LAYER Metal2 ;
        RECT 372.425 109.960 372.735 109.990 ;
        RECT 372.425 103.860 372.740 109.960 ;
        RECT 385.925 101.865 386.255 112.560 ;
    END
  END b3_c3
  PIN b4_c0_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 558.025 171.230 559.480 171.610 ;
        RECT 558.185 168.930 559.480 169.310 ;
        RECT 571.670 168.930 572.980 169.310 ;
        RECT 556.515 167.605 572.525 167.980 ;
        RECT 558.195 163.430 559.500 163.810 ;
        RECT 571.535 163.430 573.000 163.810 ;
        RECT 558.010 161.430 559.500 161.810 ;
      LAYER Metal2 ;
        RECT 558.315 160.720 558.670 171.805 ;
        RECT 571.825 163.150 572.155 169.345 ;
    END
  END b4_c0_not
  PIN b4_c1_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 557.940 151.515 559.395 151.895 ;
        RECT 558.100 149.215 559.395 149.595 ;
        RECT 571.585 149.215 572.895 149.595 ;
        RECT 556.430 147.890 572.440 148.265 ;
        RECT 558.110 143.715 559.415 144.095 ;
        RECT 571.450 143.715 572.915 144.095 ;
        RECT 557.925 141.715 559.415 142.095 ;
      LAYER Metal2 ;
        RECT 558.230 141.005 558.585 152.090 ;
        RECT 571.740 143.435 572.070 149.630 ;
    END
  END b4_c1_not
  PIN b4_c0
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 581.720 171.330 583.000 171.710 ;
        RECT 568.220 168.930 569.405 169.310 ;
        RECT 581.720 168.930 582.735 169.310 ;
        RECT 556.515 166.250 582.745 166.640 ;
        RECT 568.200 163.430 569.560 163.810 ;
        RECT 581.700 163.430 582.880 163.810 ;
        RECT 581.700 161.430 582.775 161.810 ;
      LAYER Metal2 ;
        RECT 568.840 169.295 569.150 169.325 ;
        RECT 568.840 163.195 569.155 169.295 ;
        RECT 582.340 161.200 582.670 171.895 ;
    END
  END b4_c0
  PIN b4_c1
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 581.635 151.615 582.915 151.995 ;
        RECT 568.135 149.215 569.320 149.595 ;
        RECT 581.635 149.215 582.650 149.595 ;
        RECT 556.430 146.535 582.660 146.925 ;
        RECT 568.115 143.715 569.475 144.095 ;
        RECT 581.615 143.715 582.795 144.095 ;
        RECT 581.615 141.715 582.690 142.095 ;
      LAYER Metal2 ;
        RECT 568.755 149.580 569.065 149.610 ;
        RECT 568.755 143.480 569.070 149.580 ;
        RECT 582.255 141.485 582.585 152.180 ;
    END
  END b4_c1
  PIN b4_c2_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 558.000 131.710 559.455 132.090 ;
        RECT 558.160 129.410 559.455 129.790 ;
        RECT 571.645 129.410 572.955 129.790 ;
        RECT 556.490 128.085 572.500 128.460 ;
        RECT 558.170 123.910 559.475 124.290 ;
        RECT 571.510 123.910 572.975 124.290 ;
        RECT 557.985 121.910 559.475 122.290 ;
      LAYER Metal2 ;
        RECT 558.290 121.200 558.645 132.285 ;
        RECT 571.800 123.630 572.130 129.825 ;
    END
  END b4_c2_not
  PIN b4_c2
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 581.695 131.810 582.975 132.190 ;
        RECT 568.195 129.410 569.380 129.790 ;
        RECT 581.695 129.410 582.710 129.790 ;
        RECT 556.490 126.730 582.720 127.120 ;
        RECT 568.175 123.910 569.535 124.290 ;
        RECT 581.675 123.910 582.855 124.290 ;
        RECT 581.675 121.910 582.750 122.290 ;
      LAYER Metal2 ;
        RECT 568.815 129.775 569.125 129.805 ;
        RECT 568.815 123.675 569.130 129.775 ;
        RECT 582.315 121.680 582.645 132.375 ;
    END
  END b4_c2
  PIN b4_c3_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 557.930 111.940 559.385 112.320 ;
        RECT 558.090 109.640 559.385 110.020 ;
        RECT 571.575 109.640 572.885 110.020 ;
        RECT 556.420 108.315 572.430 108.690 ;
        RECT 558.100 104.140 559.405 104.520 ;
        RECT 571.440 104.140 572.905 104.520 ;
        RECT 557.915 102.140 559.405 102.520 ;
      LAYER Metal2 ;
        RECT 558.220 101.430 558.575 112.515 ;
        RECT 571.730 103.860 572.060 110.055 ;
    END
  END b4_c3_not
  PIN b4_c3
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 581.625 112.040 582.905 112.420 ;
        RECT 568.125 109.640 569.310 110.020 ;
        RECT 581.625 109.640 582.640 110.020 ;
        RECT 556.420 106.960 582.650 107.350 ;
        RECT 568.105 104.140 569.465 104.520 ;
        RECT 581.605 104.140 582.785 104.520 ;
        RECT 581.605 102.140 582.680 102.520 ;
      LAYER Metal2 ;
        RECT 568.745 110.005 569.055 110.035 ;
        RECT 568.745 103.905 569.060 110.005 ;
        RECT 582.245 101.910 582.575 112.605 ;
    END
  END b4_c3
  PIN b2_q0
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT 142.075 204.210 143.695 204.535 ;
        RECT 166.950 168.225 167.330 168.605 ;
        RECT 188.450 168.225 188.830 168.605 ;
        RECT 163.805 165.880 182.475 165.890 ;
        RECT 142.890 165.570 190.460 165.880 ;
        RECT 142.890 165.555 164.100 165.570 ;
        RECT 174.950 163.110 175.330 163.115 ;
        RECT 172.470 162.745 175.335 163.110 ;
        RECT 180.450 163.090 180.830 163.115 ;
        RECT 180.435 162.770 182.580 163.090 ;
        RECT 174.950 162.735 175.330 162.745 ;
        RECT 180.450 162.735 180.830 162.770 ;
        RECT 166.865 148.510 167.245 148.890 ;
        RECT 188.365 148.510 188.745 148.890 ;
        RECT 142.910 146.175 163.930 146.185 ;
        RECT 142.910 146.165 182.390 146.175 ;
        RECT 142.910 145.860 190.375 146.165 ;
        RECT 163.720 145.855 190.375 145.860 ;
        RECT 174.865 143.395 175.245 143.400 ;
        RECT 172.385 143.030 175.250 143.395 ;
        RECT 180.365 143.375 180.745 143.400 ;
        RECT 180.350 143.055 182.495 143.375 ;
        RECT 174.865 143.020 175.245 143.030 ;
        RECT 180.365 143.020 180.745 143.055 ;
        RECT 166.925 128.705 167.305 129.085 ;
        RECT 188.425 128.705 188.805 129.085 ;
        RECT 142.860 126.370 164.140 126.375 ;
        RECT 142.860 126.360 182.450 126.370 ;
        RECT 142.860 126.050 190.435 126.360 ;
        RECT 174.925 123.590 175.305 123.595 ;
        RECT 172.445 123.225 175.310 123.590 ;
        RECT 180.425 123.570 180.805 123.595 ;
        RECT 180.410 123.250 182.555 123.570 ;
        RECT 174.925 123.215 175.305 123.225 ;
        RECT 180.425 123.215 180.805 123.250 ;
        RECT 166.855 108.935 167.235 109.315 ;
        RECT 188.355 108.935 188.735 109.315 ;
        RECT 142.865 106.600 163.910 106.615 ;
        RECT 142.865 106.590 182.380 106.600 ;
        RECT 142.865 106.290 190.365 106.590 ;
        RECT 163.710 106.280 190.365 106.290 ;
        RECT 174.855 103.820 175.235 103.825 ;
        RECT 172.375 103.455 175.240 103.820 ;
        RECT 180.355 103.800 180.735 103.825 ;
        RECT 180.340 103.480 182.485 103.800 ;
        RECT 174.855 103.445 175.235 103.455 ;
        RECT 180.355 103.445 180.735 103.480 ;
        RECT 166.885 89.210 167.265 89.590 ;
        RECT 188.385 89.210 188.765 89.590 ;
        RECT 142.850 86.875 163.930 86.880 ;
        RECT 142.850 86.865 182.410 86.875 ;
        RECT 142.850 86.555 190.395 86.865 ;
        RECT 174.885 84.095 175.265 84.100 ;
        RECT 172.405 83.730 175.270 84.095 ;
        RECT 180.385 84.075 180.765 84.100 ;
        RECT 180.370 83.755 182.515 84.075 ;
        RECT 174.885 83.720 175.265 83.730 ;
        RECT 180.385 83.720 180.765 83.755 ;
        RECT 166.815 69.380 167.195 69.760 ;
        RECT 188.315 69.380 188.695 69.760 ;
        RECT 142.835 67.035 182.340 67.045 ;
        RECT 142.835 66.725 190.325 67.035 ;
        RECT 142.835 66.720 163.855 66.725 ;
        RECT 174.815 64.265 175.195 64.270 ;
        RECT 172.335 63.900 175.200 64.265 ;
        RECT 180.315 64.245 180.695 64.270 ;
        RECT 180.300 63.925 182.445 64.245 ;
        RECT 174.815 63.890 175.195 63.900 ;
        RECT 180.315 63.890 180.695 63.925 ;
        RECT 166.885 49.660 167.265 50.040 ;
        RECT 188.385 49.660 188.765 50.040 ;
        RECT 142.945 47.325 163.995 47.335 ;
        RECT 142.945 47.315 182.410 47.325 ;
        RECT 142.945 47.010 190.395 47.315 ;
        RECT 163.740 47.005 190.395 47.010 ;
        RECT 174.885 44.545 175.265 44.550 ;
        RECT 172.405 44.180 175.270 44.545 ;
        RECT 180.385 44.525 180.765 44.550 ;
        RECT 180.370 44.205 182.515 44.525 ;
        RECT 174.885 44.170 175.265 44.180 ;
        RECT 180.385 44.170 180.765 44.205 ;
        RECT 166.860 29.930 167.240 30.310 ;
        RECT 188.360 29.930 188.740 30.310 ;
        RECT 163.715 27.590 182.385 27.595 ;
        RECT 142.880 27.585 182.385 27.590 ;
        RECT 142.880 27.275 190.370 27.585 ;
        RECT 142.880 27.265 163.860 27.275 ;
        RECT 174.860 24.815 175.240 24.820 ;
        RECT 172.380 24.450 175.245 24.815 ;
        RECT 180.360 24.795 180.740 24.820 ;
        RECT 180.345 24.475 182.490 24.795 ;
        RECT 174.860 24.440 175.240 24.450 ;
        RECT 180.360 24.440 180.740 24.475 ;
      LAYER Metal2 ;
        RECT 143.100 17.840 143.495 204.535 ;
        RECT 166.900 165.570 167.350 168.560 ;
        RECT 172.625 162.560 173.030 165.890 ;
        RECT 182.060 162.615 182.510 165.890 ;
        RECT 188.415 165.570 188.865 168.580 ;
        RECT 166.815 145.855 167.265 148.845 ;
        RECT 172.540 142.845 172.945 146.175 ;
        RECT 181.975 142.900 182.425 146.175 ;
        RECT 188.330 145.855 188.780 148.865 ;
        RECT 166.875 126.050 167.325 129.040 ;
        RECT 172.600 123.040 173.005 126.370 ;
        RECT 182.035 123.095 182.485 126.370 ;
        RECT 188.390 126.050 188.840 129.060 ;
        RECT 166.805 106.280 167.255 109.270 ;
        RECT 172.530 103.270 172.935 106.600 ;
        RECT 181.965 103.325 182.415 106.600 ;
        RECT 188.320 106.280 188.770 109.290 ;
        RECT 166.835 86.555 167.285 89.545 ;
        RECT 172.560 83.545 172.965 86.875 ;
        RECT 181.995 83.600 182.445 86.875 ;
        RECT 188.350 86.555 188.800 89.565 ;
        RECT 166.765 66.725 167.215 69.715 ;
        RECT 172.490 63.715 172.895 67.045 ;
        RECT 181.925 63.770 182.375 67.045 ;
        RECT 188.280 66.725 188.730 69.735 ;
        RECT 166.835 47.005 167.285 49.995 ;
        RECT 172.560 43.995 172.965 47.325 ;
        RECT 181.995 44.050 182.445 47.325 ;
        RECT 188.350 47.005 188.800 50.015 ;
        RECT 166.810 27.275 167.260 30.265 ;
        RECT 172.535 24.265 172.940 27.595 ;
        RECT 181.970 24.320 182.420 27.595 ;
        RECT 188.325 27.275 188.775 30.285 ;
    END
  END b2_q0
  PIN b2_q0_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT 142.060 203.635 144.620 203.940 ;
        RECT 170.950 168.225 171.330 168.605 ;
        RECT 184.450 168.225 184.830 168.605 ;
        RECT 163.805 164.890 190.460 164.900 ;
        RECT 144.050 164.630 190.460 164.890 ;
        RECT 144.050 164.620 164.045 164.630 ;
        RECT 166.950 163.080 167.330 163.115 ;
        RECT 188.450 163.095 188.830 163.115 ;
        RECT 166.685 162.770 169.695 163.080 ;
        RECT 185.985 162.775 188.895 163.095 ;
        RECT 166.950 162.735 167.330 162.770 ;
        RECT 188.450 162.735 188.830 162.775 ;
        RECT 170.865 148.510 171.245 148.890 ;
        RECT 184.365 148.510 184.745 148.890 ;
        RECT 144.070 145.185 163.875 145.195 ;
        RECT 144.070 144.925 190.375 145.185 ;
        RECT 163.720 144.915 190.375 144.925 ;
        RECT 166.865 143.365 167.245 143.400 ;
        RECT 188.365 143.380 188.745 143.400 ;
        RECT 166.600 143.055 169.610 143.365 ;
        RECT 185.900 143.060 188.810 143.380 ;
        RECT 166.865 143.020 167.245 143.055 ;
        RECT 188.365 143.020 188.745 143.060 ;
        RECT 170.925 128.705 171.305 129.085 ;
        RECT 184.425 128.705 184.805 129.085 ;
        RECT 144.020 125.380 164.105 125.385 ;
        RECT 144.020 125.115 190.435 125.380 ;
        RECT 163.780 125.110 190.435 125.115 ;
        RECT 166.925 123.560 167.305 123.595 ;
        RECT 188.425 123.575 188.805 123.595 ;
        RECT 166.660 123.250 169.670 123.560 ;
        RECT 185.960 123.255 188.870 123.575 ;
        RECT 166.925 123.215 167.305 123.250 ;
        RECT 188.425 123.215 188.805 123.255 ;
        RECT 170.855 108.935 171.235 109.315 ;
        RECT 184.355 108.935 184.735 109.315 ;
        RECT 144.025 105.610 163.930 105.625 ;
        RECT 144.025 105.355 190.365 105.610 ;
        RECT 163.710 105.340 190.365 105.355 ;
        RECT 166.855 103.790 167.235 103.825 ;
        RECT 188.355 103.805 188.735 103.825 ;
        RECT 166.590 103.480 169.600 103.790 ;
        RECT 185.890 103.485 188.800 103.805 ;
        RECT 166.855 103.445 167.235 103.480 ;
        RECT 188.355 103.445 188.735 103.485 ;
        RECT 170.885 89.210 171.265 89.590 ;
        RECT 184.385 89.210 184.765 89.590 ;
        RECT 144.010 85.885 163.985 85.890 ;
        RECT 144.010 85.620 190.395 85.885 ;
        RECT 163.740 85.615 190.395 85.620 ;
        RECT 166.885 84.065 167.265 84.100 ;
        RECT 188.385 84.080 188.765 84.100 ;
        RECT 166.620 83.755 169.630 84.065 ;
        RECT 185.920 83.760 188.830 84.080 ;
        RECT 166.885 83.720 167.265 83.755 ;
        RECT 188.385 83.720 188.765 83.760 ;
        RECT 170.815 69.380 171.195 69.760 ;
        RECT 184.315 69.380 184.695 69.760 ;
        RECT 143.990 65.785 190.325 66.055 ;
        RECT 166.815 64.235 167.195 64.270 ;
        RECT 188.315 64.250 188.695 64.270 ;
        RECT 166.550 63.925 169.560 64.235 ;
        RECT 185.850 63.930 188.760 64.250 ;
        RECT 166.815 63.890 167.195 63.925 ;
        RECT 188.315 63.890 188.695 63.930 ;
        RECT 170.885 49.660 171.265 50.040 ;
        RECT 184.385 49.660 184.765 50.040 ;
        RECT 144.105 46.335 163.995 46.345 ;
        RECT 144.105 46.075 190.395 46.335 ;
        RECT 163.740 46.065 190.395 46.075 ;
        RECT 166.885 44.515 167.265 44.550 ;
        RECT 188.385 44.530 188.765 44.550 ;
        RECT 166.620 44.205 169.630 44.515 ;
        RECT 185.920 44.210 188.830 44.530 ;
        RECT 166.885 44.170 167.265 44.205 ;
        RECT 188.385 44.170 188.765 44.210 ;
        RECT 170.860 29.930 171.240 30.310 ;
        RECT 184.360 29.930 184.740 30.310 ;
        RECT 163.715 26.600 190.370 26.605 ;
        RECT 144.040 26.335 190.370 26.600 ;
        RECT 144.040 26.330 163.940 26.335 ;
        RECT 166.860 24.785 167.240 24.820 ;
        RECT 188.360 24.800 188.740 24.820 ;
        RECT 166.595 24.475 169.605 24.785 ;
        RECT 185.895 24.480 188.805 24.800 ;
        RECT 166.860 24.440 167.240 24.475 ;
        RECT 188.360 24.440 188.740 24.480 ;
      LAYER Metal2 ;
        RECT 144.205 17.925 144.545 204.525 ;
        RECT 169.300 162.585 169.595 164.955 ;
        RECT 170.910 164.630 171.360 168.595 ;
        RECT 184.440 164.630 184.840 168.570 ;
        RECT 186.090 162.620 186.505 165.010 ;
        RECT 169.215 142.870 169.510 145.240 ;
        RECT 170.825 144.915 171.275 148.880 ;
        RECT 184.355 144.915 184.755 148.855 ;
        RECT 186.005 142.905 186.420 145.295 ;
        RECT 169.275 123.065 169.570 125.435 ;
        RECT 170.885 125.110 171.335 129.075 ;
        RECT 184.415 125.110 184.815 129.050 ;
        RECT 186.065 123.100 186.480 125.490 ;
        RECT 169.205 103.295 169.500 105.665 ;
        RECT 170.815 105.340 171.265 109.305 ;
        RECT 184.345 105.340 184.745 109.280 ;
        RECT 185.995 103.330 186.410 105.720 ;
        RECT 169.235 83.570 169.530 85.940 ;
        RECT 170.845 85.615 171.295 89.580 ;
        RECT 184.375 85.615 184.775 89.555 ;
        RECT 186.025 83.605 186.440 85.995 ;
        RECT 169.165 63.740 169.460 66.110 ;
        RECT 170.775 65.785 171.225 69.750 ;
        RECT 184.305 65.785 184.705 69.725 ;
        RECT 185.955 63.775 186.370 66.165 ;
        RECT 169.235 44.020 169.530 46.390 ;
        RECT 170.845 46.065 171.295 50.030 ;
        RECT 184.375 46.065 184.775 50.005 ;
        RECT 186.025 44.055 186.440 46.445 ;
        RECT 169.210 24.290 169.505 26.660 ;
        RECT 170.820 26.335 171.270 30.300 ;
        RECT 184.350 26.335 184.750 30.275 ;
        RECT 186.000 24.325 186.415 26.715 ;
    END
  END b2_q0_not
  PIN b2_c0_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 165.315 171.225 166.770 171.605 ;
        RECT 165.475 168.925 166.770 169.305 ;
        RECT 178.960 168.925 180.270 169.305 ;
        RECT 163.805 167.600 179.815 167.975 ;
        RECT 165.485 163.425 166.790 163.805 ;
        RECT 178.825 163.425 180.290 163.805 ;
        RECT 165.300 161.425 166.790 161.805 ;
      LAYER Metal2 ;
        RECT 165.605 160.715 165.960 171.800 ;
        RECT 179.115 163.145 179.445 169.340 ;
    END
  END b2_c0_not
  PIN b2_c0
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 189.010 171.325 190.290 171.705 ;
        RECT 175.510 168.925 176.695 169.305 ;
        RECT 189.010 168.925 190.025 169.305 ;
        RECT 163.805 166.245 190.035 166.635 ;
        RECT 175.490 163.425 176.850 163.805 ;
        RECT 188.990 163.425 190.170 163.805 ;
        RECT 188.990 161.425 190.065 161.805 ;
      LAYER Metal2 ;
        RECT 176.130 169.290 176.440 169.320 ;
        RECT 176.130 163.190 176.445 169.290 ;
        RECT 189.630 161.195 189.960 171.890 ;
    END
  END b2_c0
  PIN x0_c0_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 107.905 168.860 108.285 169.240 ;
        RECT 105.230 168.435 106.970 168.725 ;
        RECT 118.435 167.675 134.355 167.975 ;
        RECT 120.165 165.020 124.295 165.320 ;
        RECT 126.670 164.970 131.170 165.280 ;
        RECT 106.585 163.840 117.065 164.175 ;
        RECT 106.555 162.520 108.335 162.810 ;
        RECT 105.285 161.905 105.665 162.285 ;
      LAYER Metal2 ;
        RECT 105.315 161.845 105.615 168.775 ;
        RECT 106.625 162.445 106.925 168.795 ;
        RECT 107.940 162.475 108.235 169.300 ;
        RECT 116.625 163.810 117.005 164.190 ;
        RECT 118.475 163.690 118.790 168.015 ;
      LAYER Metal3 ;
        RECT 116.580 163.790 118.865 164.215 ;
    END
  END x0_c0_b
  PIN x0_c0_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 114.805 168.850 115.185 169.230 ;
        RECT 111.730 168.345 114.360 168.800 ;
        RECT 118.970 166.930 135.915 167.230 ;
        RECT 113.915 165.915 117.045 166.190 ;
        RECT 121.395 163.255 124.315 163.555 ;
        RECT 127.860 163.240 131.230 163.540 ;
        RECT 113.930 162.490 115.240 162.810 ;
        RECT 111.740 161.935 112.120 162.315 ;
      LAYER Metal2 ;
        RECT 111.780 161.845 112.080 168.785 ;
        RECT 113.990 162.420 114.270 168.780 ;
        RECT 114.840 162.420 115.140 169.240 ;
        RECT 116.625 165.865 117.005 166.245 ;
        RECT 119.085 165.765 119.365 167.295 ;
        RECT 121.430 163.205 121.730 167.265 ;
        RECT 127.920 163.190 128.200 167.280 ;
      LAYER Metal3 ;
        RECT 116.605 165.865 119.450 166.245 ;
    END
  END x0_c0_b_not
  PIN p1
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 123.365 168.860 123.745 169.240 ;
        RECT 120.690 168.435 122.430 168.725 ;
        RECT 122.045 163.840 138.065 164.175 ;
        RECT 122.015 162.520 123.795 162.810 ;
        RECT 120.745 161.905 121.125 162.285 ;
      LAYER Metal2 ;
        RECT 120.775 161.845 121.075 168.775 ;
        RECT 122.085 162.445 122.385 168.795 ;
        RECT 123.400 162.475 123.695 169.300 ;
    END
  END p1
  PIN p1_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 130.265 168.850 130.645 169.230 ;
        RECT 127.190 168.355 129.815 168.765 ;
        RECT 129.375 165.915 137.075 166.190 ;
        RECT 129.390 162.490 130.700 162.810 ;
        RECT 127.200 161.935 127.580 162.315 ;
      LAYER Metal2 ;
        RECT 127.240 161.845 127.540 168.785 ;
        RECT 129.450 162.420 129.730 168.780 ;
        RECT 130.300 162.420 130.600 169.240 ;
    END
  END p1_not
  PIN b0_q1
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -54.095 204.200 -52.475 204.525 ;
        RECT -29.310 187.870 -28.930 188.250 ;
        RECT -7.810 187.870 -7.430 188.250 ;
        RECT -53.285 185.535 -32.075 185.620 ;
        RECT -53.285 185.525 -13.785 185.535 ;
        RECT -53.285 185.295 -5.800 185.525 ;
        RECT -32.455 185.215 -5.800 185.295 ;
        RECT -21.310 182.755 -20.930 182.760 ;
        RECT -23.790 182.390 -20.925 182.755 ;
        RECT -15.810 182.735 -15.430 182.760 ;
        RECT -15.825 182.415 -13.680 182.735 ;
        RECT -21.310 182.380 -20.930 182.390 ;
        RECT -15.810 182.380 -15.430 182.415 ;
        RECT -29.220 168.215 -28.840 168.595 ;
        RECT -7.720 168.215 -7.340 168.595 ;
        RECT -53.250 165.880 -32.230 165.905 ;
        RECT -53.250 165.870 -13.695 165.880 ;
        RECT -53.250 165.580 -5.710 165.870 ;
        RECT -32.365 165.560 -5.710 165.580 ;
        RECT -21.220 163.100 -20.840 163.105 ;
        RECT -23.700 162.735 -20.835 163.100 ;
        RECT -15.720 163.080 -15.340 163.105 ;
        RECT -15.735 162.760 -13.590 163.080 ;
        RECT -21.220 162.725 -20.840 162.735 ;
        RECT -15.720 162.725 -15.340 162.760 ;
        RECT -29.305 148.500 -28.925 148.880 ;
        RECT -7.805 148.500 -7.425 148.880 ;
        RECT -32.450 146.155 -13.780 146.165 ;
        RECT -32.450 146.095 -5.795 146.155 ;
        RECT -53.300 145.845 -5.795 146.095 ;
        RECT -53.300 145.770 -32.020 145.845 ;
        RECT -21.305 143.385 -20.925 143.390 ;
        RECT -23.785 143.020 -20.920 143.385 ;
        RECT -15.805 143.365 -15.425 143.390 ;
        RECT -15.820 143.045 -13.675 143.365 ;
        RECT -21.305 143.010 -20.925 143.020 ;
        RECT -15.805 143.010 -15.425 143.045 ;
        RECT -29.245 128.695 -28.865 129.075 ;
        RECT -7.745 128.695 -7.365 129.075 ;
        RECT -32.390 126.350 -13.720 126.360 ;
        RECT -32.390 126.335 -5.735 126.350 ;
        RECT -53.295 126.040 -5.735 126.335 ;
        RECT -53.295 126.010 -32.250 126.040 ;
        RECT -21.245 123.580 -20.865 123.585 ;
        RECT -23.725 123.215 -20.860 123.580 ;
        RECT -15.745 123.560 -15.365 123.585 ;
        RECT -15.760 123.240 -13.615 123.560 ;
        RECT -21.245 123.205 -20.865 123.215 ;
        RECT -15.745 123.205 -15.365 123.240 ;
        RECT -29.315 108.925 -28.935 109.305 ;
        RECT -7.815 108.925 -7.435 109.305 ;
        RECT -53.310 106.590 -32.230 106.600 ;
        RECT -53.310 106.580 -13.790 106.590 ;
        RECT -53.310 106.275 -5.805 106.580 ;
        RECT -32.460 106.270 -5.805 106.275 ;
        RECT -21.315 103.810 -20.935 103.815 ;
        RECT -23.795 103.445 -20.930 103.810 ;
        RECT -15.815 103.790 -15.435 103.815 ;
        RECT -15.830 103.470 -13.685 103.790 ;
        RECT -21.315 103.435 -20.935 103.445 ;
        RECT -15.815 103.435 -15.435 103.470 ;
        RECT -29.285 89.200 -28.905 89.580 ;
        RECT -7.785 89.200 -7.405 89.580 ;
        RECT -32.430 86.860 -13.760 86.865 ;
        RECT -53.330 86.855 -13.760 86.860 ;
        RECT -53.330 86.545 -5.775 86.855 ;
        RECT -53.330 86.535 -32.310 86.545 ;
        RECT -21.285 84.085 -20.905 84.090 ;
        RECT -23.765 83.720 -20.900 84.085 ;
        RECT -15.785 84.065 -15.405 84.090 ;
        RECT -15.800 83.745 -13.655 84.065 ;
        RECT -21.285 83.710 -20.905 83.720 ;
        RECT -15.785 83.710 -15.405 83.745 ;
        RECT -29.355 69.370 -28.975 69.750 ;
        RECT -7.855 69.370 -7.475 69.750 ;
        RECT -53.215 67.035 -32.165 67.055 ;
        RECT -53.215 67.025 -13.830 67.035 ;
        RECT -53.215 66.730 -5.845 67.025 ;
        RECT -32.500 66.715 -5.845 66.730 ;
        RECT -21.355 64.255 -20.975 64.260 ;
        RECT -23.835 63.890 -20.970 64.255 ;
        RECT -15.855 64.235 -15.475 64.260 ;
        RECT -15.870 63.915 -13.725 64.235 ;
        RECT -21.355 63.880 -20.975 63.890 ;
        RECT -15.855 63.880 -15.475 63.915 ;
        RECT -29.285 49.650 -28.905 50.030 ;
        RECT -7.785 49.650 -7.405 50.030 ;
        RECT -32.430 47.310 -13.760 47.315 ;
        RECT -53.280 47.305 -13.760 47.310 ;
        RECT -53.280 46.995 -5.775 47.305 ;
        RECT -53.280 46.985 -32.300 46.995 ;
        RECT -21.285 44.535 -20.905 44.540 ;
        RECT -23.765 44.170 -20.900 44.535 ;
        RECT -15.785 44.515 -15.405 44.540 ;
        RECT -15.800 44.195 -13.655 44.515 ;
        RECT -21.285 44.160 -20.905 44.170 ;
        RECT -15.785 44.160 -15.405 44.195 ;
      LAYER Metal2 ;
        RECT -53.070 17.830 -52.675 204.525 ;
        RECT -29.360 185.215 -28.910 188.205 ;
        RECT -23.635 182.205 -23.230 185.535 ;
        RECT -14.200 182.260 -13.750 185.535 ;
        RECT -7.845 185.215 -7.395 188.225 ;
        RECT -29.270 165.560 -28.820 168.550 ;
        RECT -23.545 162.550 -23.140 165.880 ;
        RECT -14.110 162.605 -13.660 165.880 ;
        RECT -7.755 165.560 -7.305 168.570 ;
        RECT -29.355 145.845 -28.905 148.835 ;
        RECT -23.630 142.835 -23.225 146.165 ;
        RECT -14.195 142.890 -13.745 146.165 ;
        RECT -7.840 145.845 -7.390 148.855 ;
        RECT -29.295 126.040 -28.845 129.030 ;
        RECT -23.570 123.030 -23.165 126.360 ;
        RECT -14.135 123.085 -13.685 126.360 ;
        RECT -7.780 126.040 -7.330 129.050 ;
        RECT -29.365 106.270 -28.915 109.260 ;
        RECT -23.640 103.260 -23.235 106.590 ;
        RECT -14.205 103.315 -13.755 106.590 ;
        RECT -7.850 106.270 -7.400 109.280 ;
        RECT -29.335 86.545 -28.885 89.535 ;
        RECT -23.610 83.535 -23.205 86.865 ;
        RECT -14.175 83.590 -13.725 86.865 ;
        RECT -7.820 86.545 -7.370 89.555 ;
        RECT -29.405 66.715 -28.955 69.705 ;
        RECT -23.680 63.705 -23.275 67.035 ;
        RECT -14.245 63.760 -13.795 67.035 ;
        RECT -7.890 66.715 -7.440 69.725 ;
        RECT -29.335 46.995 -28.885 49.985 ;
        RECT -23.610 43.985 -23.205 47.315 ;
        RECT -14.175 44.040 -13.725 47.315 ;
        RECT -7.820 46.995 -7.370 50.005 ;
    END
  END b0_q1
  PIN b0_q1_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -54.110 203.625 -51.550 203.930 ;
        RECT -25.310 187.870 -24.930 188.250 ;
        RECT -11.810 187.870 -11.430 188.250 ;
        RECT -52.125 184.545 -32.130 184.630 ;
        RECT -52.125 184.360 -5.800 184.545 ;
        RECT -32.455 184.275 -5.800 184.360 ;
        RECT -29.310 182.725 -28.930 182.760 ;
        RECT -7.810 182.740 -7.430 182.760 ;
        RECT -29.575 182.415 -26.565 182.725 ;
        RECT -10.275 182.420 -7.365 182.740 ;
        RECT -29.310 182.380 -28.930 182.415 ;
        RECT -7.810 182.380 -7.430 182.420 ;
        RECT -25.220 168.215 -24.840 168.595 ;
        RECT -11.720 168.215 -11.340 168.595 ;
        RECT -52.090 164.890 -32.285 164.915 ;
        RECT -52.090 164.645 -5.710 164.890 ;
        RECT -32.365 164.620 -5.710 164.645 ;
        RECT -29.220 163.070 -28.840 163.105 ;
        RECT -7.720 163.085 -7.340 163.105 ;
        RECT -29.485 162.760 -26.475 163.070 ;
        RECT -10.185 162.765 -7.275 163.085 ;
        RECT -29.220 162.725 -28.840 162.760 ;
        RECT -7.720 162.725 -7.340 162.765 ;
        RECT -25.305 148.500 -24.925 148.880 ;
        RECT -11.805 148.500 -11.425 148.880 ;
        RECT -32.450 145.105 -5.795 145.175 ;
        RECT -52.140 144.905 -5.795 145.105 ;
        RECT -52.140 144.835 -32.055 144.905 ;
        RECT -29.305 143.355 -28.925 143.390 ;
        RECT -7.805 143.370 -7.425 143.390 ;
        RECT -29.570 143.045 -26.560 143.355 ;
        RECT -10.270 143.050 -7.360 143.370 ;
        RECT -29.305 143.010 -28.925 143.045 ;
        RECT -7.805 143.010 -7.425 143.050 ;
        RECT -25.245 128.695 -24.865 129.075 ;
        RECT -11.745 128.695 -11.365 129.075 ;
        RECT -32.390 125.345 -5.735 125.370 ;
        RECT -52.135 125.100 -5.735 125.345 ;
        RECT -52.135 125.075 -32.230 125.100 ;
        RECT -29.245 123.550 -28.865 123.585 ;
        RECT -7.745 123.565 -7.365 123.585 ;
        RECT -29.510 123.240 -26.500 123.550 ;
        RECT -10.210 123.245 -7.300 123.565 ;
        RECT -29.245 123.205 -28.865 123.240 ;
        RECT -7.745 123.205 -7.365 123.245 ;
        RECT -25.315 108.925 -24.935 109.305 ;
        RECT -11.815 108.925 -11.435 109.305 ;
        RECT -52.150 105.600 -32.175 105.610 ;
        RECT -52.150 105.340 -5.805 105.600 ;
        RECT -32.460 105.330 -5.805 105.340 ;
        RECT -29.315 103.780 -28.935 103.815 ;
        RECT -7.815 103.795 -7.435 103.815 ;
        RECT -29.580 103.470 -26.570 103.780 ;
        RECT -10.280 103.475 -7.370 103.795 ;
        RECT -29.315 103.435 -28.935 103.470 ;
        RECT -7.815 103.435 -7.435 103.475 ;
        RECT -25.285 89.200 -24.905 89.580 ;
        RECT -11.785 89.200 -11.405 89.580 ;
        RECT -32.430 85.870 -5.775 85.875 ;
        RECT -52.170 85.605 -5.775 85.870 ;
        RECT -52.170 85.600 -32.370 85.605 ;
        RECT -29.285 84.055 -28.905 84.090 ;
        RECT -7.785 84.070 -7.405 84.090 ;
        RECT -29.550 83.745 -26.540 84.055 ;
        RECT -10.250 83.750 -7.340 84.070 ;
        RECT -29.285 83.710 -28.905 83.745 ;
        RECT -7.785 83.710 -7.405 83.750 ;
        RECT -25.355 69.370 -24.975 69.750 ;
        RECT -11.855 69.370 -11.475 69.750 ;
        RECT -52.055 66.045 -32.165 66.065 ;
        RECT -52.055 65.795 -5.845 66.045 ;
        RECT -32.500 65.775 -5.845 65.795 ;
        RECT -29.355 64.225 -28.975 64.260 ;
        RECT -7.855 64.240 -7.475 64.260 ;
        RECT -29.620 63.915 -26.610 64.225 ;
        RECT -10.320 63.920 -7.410 64.240 ;
        RECT -29.355 63.880 -28.975 63.915 ;
        RECT -7.855 63.880 -7.475 63.920 ;
        RECT -25.285 49.650 -24.905 50.030 ;
        RECT -11.785 49.650 -11.405 50.030 ;
        RECT -32.430 46.320 -5.775 46.325 ;
        RECT -52.120 46.055 -5.775 46.320 ;
        RECT -52.120 46.050 -32.220 46.055 ;
        RECT -29.285 44.505 -28.905 44.540 ;
        RECT -7.785 44.520 -7.405 44.540 ;
        RECT -29.550 44.195 -26.540 44.505 ;
        RECT -10.250 44.200 -7.340 44.520 ;
        RECT -29.285 44.160 -28.905 44.195 ;
        RECT -7.785 44.160 -7.405 44.200 ;
      LAYER Metal2 ;
        RECT -51.965 17.915 -51.625 204.515 ;
        RECT -26.960 182.230 -26.665 184.600 ;
        RECT -25.350 184.275 -24.900 188.240 ;
        RECT -11.820 184.275 -11.420 188.215 ;
        RECT -10.170 182.265 -9.755 184.655 ;
        RECT -26.870 162.575 -26.575 164.945 ;
        RECT -25.260 164.620 -24.810 168.585 ;
        RECT -11.730 164.620 -11.330 168.560 ;
        RECT -10.080 162.610 -9.665 165.000 ;
        RECT -26.955 142.860 -26.660 145.230 ;
        RECT -25.345 144.905 -24.895 148.870 ;
        RECT -11.815 144.905 -11.415 148.845 ;
        RECT -10.165 142.895 -9.750 145.285 ;
        RECT -26.895 123.055 -26.600 125.425 ;
        RECT -25.285 125.100 -24.835 129.065 ;
        RECT -11.755 125.100 -11.355 129.040 ;
        RECT -10.105 123.090 -9.690 125.480 ;
        RECT -26.965 103.285 -26.670 105.655 ;
        RECT -25.355 105.330 -24.905 109.295 ;
        RECT -11.825 105.330 -11.425 109.270 ;
        RECT -10.175 103.320 -9.760 105.710 ;
        RECT -26.935 83.560 -26.640 85.930 ;
        RECT -25.325 85.605 -24.875 89.570 ;
        RECT -11.795 85.605 -11.395 89.545 ;
        RECT -10.145 83.595 -9.730 85.985 ;
        RECT -27.005 63.730 -26.710 66.100 ;
        RECT -25.395 65.775 -24.945 69.740 ;
        RECT -11.865 65.775 -11.465 69.715 ;
        RECT -10.215 63.765 -9.800 66.155 ;
        RECT -26.935 44.010 -26.640 46.380 ;
        RECT -25.325 46.055 -24.875 50.020 ;
        RECT -11.795 46.055 -11.395 49.995 ;
        RECT -10.145 44.045 -9.730 46.435 ;
    END
  END b0_q1_not
  PIN b1_q0_not
    ANTENNAGATEAREA 3.763200 ;
    PORT
      LAYER Metal1 ;
        RECT -106.705 203.605 -101.190 203.935 ;
        RECT -75.545 168.135 -75.165 168.515 ;
        RECT -62.045 168.135 -61.665 168.515 ;
        RECT -101.890 164.540 -56.035 164.810 ;
        RECT -79.545 162.990 -79.165 163.025 ;
        RECT -58.045 163.005 -57.665 163.025 ;
        RECT -79.810 162.680 -76.800 162.990 ;
        RECT -60.510 162.685 -57.600 163.005 ;
        RECT -79.545 162.645 -79.165 162.680 ;
        RECT -58.045 162.645 -57.665 162.685 ;
        RECT -75.630 148.420 -75.250 148.800 ;
        RECT -62.130 148.420 -61.750 148.800 ;
        RECT -101.855 144.825 -56.120 145.095 ;
        RECT -79.630 143.275 -79.250 143.310 ;
        RECT -58.130 143.290 -57.750 143.310 ;
        RECT -79.895 142.965 -76.885 143.275 ;
        RECT -60.595 142.970 -57.685 143.290 ;
        RECT -79.630 142.930 -79.250 142.965 ;
        RECT -58.130 142.930 -57.750 142.970 ;
        RECT -75.570 128.615 -75.190 128.995 ;
        RECT -62.070 128.615 -61.690 128.995 ;
        RECT -82.715 125.285 -56.060 125.290 ;
        RECT -101.905 125.020 -56.060 125.285 ;
        RECT -101.905 125.015 -82.315 125.020 ;
        RECT -79.570 123.470 -79.190 123.505 ;
        RECT -58.070 123.485 -57.690 123.505 ;
        RECT -79.835 123.160 -76.825 123.470 ;
        RECT -60.535 123.165 -57.625 123.485 ;
        RECT -79.570 123.125 -79.190 123.160 ;
        RECT -58.070 123.125 -57.690 123.165 ;
        RECT -75.640 108.845 -75.260 109.225 ;
        RECT -62.140 108.845 -61.760 109.225 ;
        RECT -101.900 105.520 -82.310 105.525 ;
        RECT -101.900 105.255 -56.130 105.520 ;
        RECT -82.785 105.250 -56.130 105.255 ;
        RECT -79.640 103.700 -79.260 103.735 ;
        RECT -58.140 103.715 -57.760 103.735 ;
        RECT -79.905 103.390 -76.895 103.700 ;
        RECT -60.605 103.395 -57.695 103.715 ;
        RECT -79.640 103.355 -79.260 103.390 ;
        RECT -58.140 103.355 -57.760 103.395 ;
        RECT -75.610 89.120 -75.230 89.500 ;
        RECT -62.110 89.120 -61.730 89.500 ;
        RECT -82.755 85.790 -56.100 85.795 ;
        RECT -101.915 85.525 -56.100 85.790 ;
        RECT -101.915 85.520 -82.325 85.525 ;
        RECT -79.610 83.975 -79.230 84.010 ;
        RECT -58.110 83.990 -57.730 84.010 ;
        RECT -79.875 83.665 -76.865 83.975 ;
        RECT -60.575 83.670 -57.665 83.990 ;
        RECT -79.610 83.630 -79.230 83.665 ;
        RECT -58.110 83.630 -57.730 83.670 ;
        RECT -75.680 69.290 -75.300 69.670 ;
        RECT -62.180 69.290 -61.800 69.670 ;
        RECT -101.935 65.965 -82.345 65.980 ;
        RECT -101.935 65.710 -56.170 65.965 ;
        RECT -82.825 65.695 -56.170 65.710 ;
        RECT -79.680 64.145 -79.300 64.180 ;
        RECT -58.180 64.160 -57.800 64.180 ;
        RECT -79.945 63.835 -76.935 64.145 ;
        RECT -60.645 63.840 -57.735 64.160 ;
        RECT -79.680 63.800 -79.300 63.835 ;
        RECT -58.180 63.800 -57.800 63.840 ;
        RECT -75.610 49.570 -75.230 49.950 ;
        RECT -62.110 49.570 -61.730 49.950 ;
        RECT -101.820 45.975 -56.100 46.245 ;
        RECT -79.610 44.425 -79.230 44.460 ;
        RECT -58.110 44.440 -57.730 44.460 ;
        RECT -79.875 44.115 -76.865 44.425 ;
        RECT -60.575 44.120 -57.665 44.440 ;
        RECT -79.610 44.080 -79.230 44.115 ;
        RECT -58.110 44.080 -57.730 44.120 ;
        RECT -75.605 29.760 -75.225 30.140 ;
        RECT -62.105 29.760 -61.725 30.140 ;
        RECT -82.750 26.430 -56.095 26.435 ;
        RECT -101.815 26.165 -56.095 26.430 ;
        RECT -101.815 26.160 -82.225 26.165 ;
        RECT -79.605 24.615 -79.225 24.650 ;
        RECT -58.105 24.630 -57.725 24.650 ;
        RECT -79.870 24.305 -76.860 24.615 ;
        RECT -60.570 24.310 -57.660 24.630 ;
        RECT -79.605 24.270 -79.225 24.305 ;
        RECT -58.105 24.270 -57.725 24.310 ;
      LAYER Metal2 ;
        RECT -101.725 18.040 -101.385 204.535 ;
        RECT -77.195 162.495 -76.900 164.865 ;
        RECT -75.585 164.540 -75.135 168.505 ;
        RECT -62.055 164.540 -61.655 168.480 ;
        RECT -60.405 162.530 -59.990 164.920 ;
        RECT -77.280 142.780 -76.985 145.150 ;
        RECT -75.670 144.825 -75.220 148.790 ;
        RECT -62.140 144.825 -61.740 148.765 ;
        RECT -60.490 142.815 -60.075 145.205 ;
        RECT -77.220 122.975 -76.925 125.345 ;
        RECT -75.610 125.020 -75.160 128.985 ;
        RECT -62.080 125.020 -61.680 128.960 ;
        RECT -60.430 123.010 -60.015 125.400 ;
        RECT -77.290 103.205 -76.995 105.575 ;
        RECT -75.680 105.250 -75.230 109.215 ;
        RECT -62.150 105.250 -61.750 109.190 ;
        RECT -60.500 103.240 -60.085 105.630 ;
        RECT -77.260 83.480 -76.965 85.850 ;
        RECT -75.650 85.525 -75.200 89.490 ;
        RECT -62.120 85.525 -61.720 89.465 ;
        RECT -60.470 83.515 -60.055 85.905 ;
        RECT -77.330 63.650 -77.035 66.020 ;
        RECT -75.720 65.695 -75.270 69.660 ;
        RECT -62.190 65.695 -61.790 69.635 ;
        RECT -60.540 63.685 -60.125 66.075 ;
        RECT -77.260 43.930 -76.965 46.300 ;
        RECT -75.650 45.975 -75.200 49.940 ;
        RECT -62.120 45.975 -61.720 49.915 ;
        RECT -60.470 43.965 -60.055 46.355 ;
        RECT -77.255 24.120 -76.960 26.490 ;
        RECT -75.645 26.165 -75.195 30.130 ;
        RECT -62.115 26.165 -61.715 30.105 ;
        RECT -60.465 24.155 -60.050 26.545 ;
    END
  END b1_q0_not
  PIN b0_c0
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -7.250 190.970 -5.970 191.350 ;
        RECT -20.750 188.570 -19.565 188.950 ;
        RECT -7.250 188.570 -6.235 188.950 ;
        RECT -32.455 185.890 -6.225 186.280 ;
        RECT -20.770 183.070 -19.410 183.450 ;
        RECT -7.270 183.070 -6.090 183.450 ;
        RECT -7.270 181.070 -6.195 181.450 ;
      LAYER Metal2 ;
        RECT -20.130 188.935 -19.820 188.965 ;
        RECT -20.130 182.835 -19.815 188.935 ;
        RECT -6.630 180.840 -6.300 191.535 ;
    END
  END b0_c0
  PIN p0_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -28.750 190.870 -27.550 191.250 ;
        RECT -28.750 188.570 -25.490 188.950 ;
        RECT -28.085 186.655 -5.800 186.995 ;
        RECT -28.770 183.070 -25.470 183.450 ;
        RECT -28.770 181.070 -27.485 181.450 ;
      LAYER Metal2 ;
        RECT -27.925 180.340 -27.610 191.390 ;
    END
  END p0_not
  PIN p0
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -9.225 190.970 -7.990 191.350 ;
        RECT -11.250 188.570 -7.990 188.950 ;
        RECT -9.365 183.710 -5.800 184.045 ;
        RECT -11.270 183.070 -7.970 183.450 ;
        RECT -9.455 181.070 -7.970 181.450 ;
      LAYER Metal2 ;
        RECT -9.140 180.825 -8.825 191.510 ;
    END
  END p0
  PIN b0_c1
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -7.160 171.315 -5.880 171.695 ;
        RECT -20.660 168.915 -19.475 169.295 ;
        RECT -7.160 168.915 -6.145 169.295 ;
        RECT -32.365 166.235 -6.135 166.625 ;
        RECT -20.680 163.415 -19.320 163.795 ;
        RECT -7.180 163.415 -6.000 163.795 ;
        RECT -7.180 161.415 -6.105 161.795 ;
      LAYER Metal2 ;
        RECT -20.040 169.280 -19.730 169.310 ;
        RECT -20.040 163.180 -19.725 169.280 ;
        RECT -6.540 161.185 -6.210 171.880 ;
    END
  END b0_c1
  PIN b0_c1_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -30.855 171.215 -29.400 171.595 ;
        RECT -30.695 168.915 -29.400 169.295 ;
        RECT -17.210 168.915 -15.900 169.295 ;
        RECT -32.365 167.590 -16.355 167.965 ;
        RECT -30.685 163.415 -29.380 163.795 ;
        RECT -17.345 163.415 -15.880 163.795 ;
        RECT -30.870 161.415 -29.380 161.795 ;
      LAYER Metal2 ;
        RECT -30.565 160.705 -30.210 171.790 ;
        RECT -17.055 163.135 -16.725 169.330 ;
    END
  END b0_c1_not
  PIN b0_c0_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -30.945 190.870 -29.490 191.250 ;
        RECT -30.785 188.570 -29.490 188.950 ;
        RECT -17.300 188.570 -15.990 188.950 ;
        RECT -32.455 187.245 -16.445 187.620 ;
        RECT -30.775 183.070 -29.470 183.450 ;
        RECT -17.435 183.070 -15.970 183.450 ;
        RECT -30.960 181.070 -29.470 181.450 ;
      LAYER Metal2 ;
        RECT -30.655 180.360 -30.300 191.445 ;
        RECT -17.145 182.790 -16.815 188.985 ;
    END
  END b0_c0_not
  PIN b1_c0_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -81.180 171.135 -79.725 171.515 ;
        RECT -81.020 168.835 -79.725 169.215 ;
        RECT -67.535 168.835 -66.225 169.215 ;
        RECT -82.690 167.510 -66.680 167.885 ;
        RECT -81.010 163.335 -79.705 163.715 ;
        RECT -67.670 163.335 -66.205 163.715 ;
        RECT -81.195 161.335 -79.705 161.715 ;
      LAYER Metal2 ;
        RECT -80.890 160.625 -80.535 171.710 ;
        RECT -67.380 163.055 -67.050 169.250 ;
    END
  END b1_c0_not
  PIN b1_c0
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -57.485 171.235 -56.205 171.615 ;
        RECT -70.985 168.835 -69.800 169.215 ;
        RECT -57.485 168.835 -56.470 169.215 ;
        RECT -82.690 166.155 -56.460 166.545 ;
        RECT -71.005 163.335 -69.645 163.715 ;
        RECT -57.505 163.335 -56.325 163.715 ;
        RECT -57.505 161.335 -56.430 161.715 ;
      LAYER Metal2 ;
        RECT -70.365 169.200 -70.055 169.230 ;
        RECT -70.365 163.100 -70.050 169.200 ;
        RECT -56.865 161.105 -56.535 171.800 ;
    END
  END b1_c0
  PIN b0_c2
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -7.245 151.600 -5.965 151.980 ;
        RECT -20.745 149.200 -19.560 149.580 ;
        RECT -7.245 149.200 -6.230 149.580 ;
        RECT -32.450 146.520 -6.220 146.910 ;
        RECT -20.765 143.700 -19.405 144.080 ;
        RECT -7.265 143.700 -6.085 144.080 ;
        RECT -7.265 141.700 -6.190 142.080 ;
      LAYER Metal2 ;
        RECT -20.125 149.565 -19.815 149.595 ;
        RECT -20.125 143.465 -19.810 149.565 ;
        RECT -6.625 141.470 -6.295 152.165 ;
    END
  END b0_c2
  PIN b0_c2_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -30.940 151.500 -29.485 151.880 ;
        RECT -30.780 149.200 -29.485 149.580 ;
        RECT -17.295 149.200 -15.985 149.580 ;
        RECT -32.450 147.875 -16.440 148.250 ;
        RECT -30.770 143.700 -29.465 144.080 ;
        RECT -17.430 143.700 -15.965 144.080 ;
        RECT -30.955 141.700 -29.465 142.080 ;
      LAYER Metal2 ;
        RECT -30.650 140.990 -30.295 152.075 ;
        RECT -17.140 143.420 -16.810 149.615 ;
    END
  END b0_c2_not
  PIN b0_c3_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -30.880 131.695 -29.425 132.075 ;
        RECT -30.720 129.395 -29.425 129.775 ;
        RECT -17.235 129.395 -15.925 129.775 ;
        RECT -32.390 128.070 -16.380 128.445 ;
        RECT -30.710 123.895 -29.405 124.275 ;
        RECT -17.370 123.895 -15.905 124.275 ;
        RECT -30.895 121.895 -29.405 122.275 ;
      LAYER Metal2 ;
        RECT -30.590 121.185 -30.235 132.270 ;
        RECT -17.080 123.615 -16.750 129.810 ;
    END
  END b0_c3_not
  PIN b0_c3
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -7.185 131.795 -5.905 132.175 ;
        RECT -20.685 129.395 -19.500 129.775 ;
        RECT -7.185 129.395 -6.170 129.775 ;
        RECT -32.390 126.715 -6.160 127.105 ;
        RECT -20.705 123.895 -19.345 124.275 ;
        RECT -7.205 123.895 -6.025 124.275 ;
        RECT -7.205 121.895 -6.130 122.275 ;
      LAYER Metal2 ;
        RECT -20.065 129.760 -19.755 129.790 ;
        RECT -20.065 123.660 -19.750 129.760 ;
        RECT -6.565 121.665 -6.235 132.360 ;
    END
  END b0_c3
  PIN b0_c4_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -30.950 111.925 -29.495 112.305 ;
        RECT -30.790 109.625 -29.495 110.005 ;
        RECT -17.305 109.625 -15.995 110.005 ;
        RECT -32.460 108.300 -16.450 108.675 ;
        RECT -30.780 104.125 -29.475 104.505 ;
        RECT -17.440 104.125 -15.975 104.505 ;
        RECT -30.965 102.125 -29.475 102.505 ;
      LAYER Metal2 ;
        RECT -30.660 101.415 -30.305 112.500 ;
        RECT -17.150 103.845 -16.820 110.040 ;
    END
  END b0_c4_not
  PIN b0_c4
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -7.255 112.025 -5.975 112.405 ;
        RECT -20.755 109.625 -19.570 110.005 ;
        RECT -7.255 109.625 -6.240 110.005 ;
        RECT -32.460 106.945 -6.230 107.335 ;
        RECT -20.775 104.125 -19.415 104.505 ;
        RECT -7.275 104.125 -6.095 104.505 ;
        RECT -7.275 102.125 -6.200 102.505 ;
      LAYER Metal2 ;
        RECT -20.135 109.990 -19.825 110.020 ;
        RECT -20.135 103.890 -19.820 109.990 ;
        RECT -6.635 101.895 -6.305 112.590 ;
    END
  END b0_c4
  PIN b1_c1_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -81.265 151.420 -79.810 151.800 ;
        RECT -81.105 149.120 -79.810 149.500 ;
        RECT -67.620 149.120 -66.310 149.500 ;
        RECT -82.775 147.795 -66.765 148.170 ;
        RECT -81.095 143.620 -79.790 144.000 ;
        RECT -67.755 143.620 -66.290 144.000 ;
        RECT -81.280 141.620 -79.790 142.000 ;
      LAYER Metal2 ;
        RECT -80.975 140.910 -80.620 151.995 ;
        RECT -67.465 143.340 -67.135 149.535 ;
    END
  END b1_c1_not
  PIN b1_c1
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -57.570 151.520 -56.290 151.900 ;
        RECT -71.070 149.120 -69.885 149.500 ;
        RECT -57.570 149.120 -56.555 149.500 ;
        RECT -82.775 146.440 -56.545 146.830 ;
        RECT -71.090 143.620 -69.730 144.000 ;
        RECT -57.590 143.620 -56.410 144.000 ;
        RECT -57.590 141.620 -56.515 142.000 ;
      LAYER Metal2 ;
        RECT -70.450 149.485 -70.140 149.515 ;
        RECT -70.450 143.385 -70.135 149.485 ;
        RECT -56.950 141.390 -56.620 152.085 ;
    END
  END b1_c1
  PIN b1_c2_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -81.205 131.615 -79.750 131.995 ;
        RECT -81.045 129.315 -79.750 129.695 ;
        RECT -67.560 129.315 -66.250 129.695 ;
        RECT -82.715 127.990 -66.705 128.365 ;
        RECT -81.035 123.815 -79.730 124.195 ;
        RECT -67.695 123.815 -66.230 124.195 ;
        RECT -81.220 121.815 -79.730 122.195 ;
      LAYER Metal2 ;
        RECT -80.915 121.105 -80.560 132.190 ;
        RECT -67.405 123.535 -67.075 129.730 ;
    END
  END b1_c2_not
  PIN b1_c2
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -57.510 131.715 -56.230 132.095 ;
        RECT -71.010 129.315 -69.825 129.695 ;
        RECT -57.510 129.315 -56.495 129.695 ;
        RECT -82.715 126.635 -56.485 127.025 ;
        RECT -71.030 123.815 -69.670 124.195 ;
        RECT -57.530 123.815 -56.350 124.195 ;
        RECT -57.530 121.815 -56.455 122.195 ;
      LAYER Metal2 ;
        RECT -70.390 129.680 -70.080 129.710 ;
        RECT -70.390 123.580 -70.075 129.680 ;
        RECT -56.890 121.585 -56.560 132.280 ;
    END
  END b1_c2
  PIN b1_c3_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -81.275 111.845 -79.820 112.225 ;
        RECT -81.115 109.545 -79.820 109.925 ;
        RECT -67.630 109.545 -66.320 109.925 ;
        RECT -82.785 108.220 -66.775 108.595 ;
        RECT -81.105 104.045 -79.800 104.425 ;
        RECT -67.765 104.045 -66.300 104.425 ;
        RECT -81.290 102.045 -79.800 102.425 ;
      LAYER Metal2 ;
        RECT -80.985 101.335 -80.630 112.420 ;
        RECT -67.475 103.765 -67.145 109.960 ;
    END
  END b1_c3_not
  PIN b1_c3
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -57.580 111.945 -56.300 112.325 ;
        RECT -71.080 109.545 -69.895 109.925 ;
        RECT -57.580 109.545 -56.565 109.925 ;
        RECT -82.785 106.865 -56.555 107.255 ;
        RECT -71.100 104.045 -69.740 104.425 ;
        RECT -57.600 104.045 -56.420 104.425 ;
        RECT -57.600 102.045 -56.525 102.425 ;
      LAYER Metal2 ;
        RECT -70.460 109.910 -70.150 109.940 ;
        RECT -70.460 103.810 -70.145 109.910 ;
        RECT -56.960 101.815 -56.630 112.510 ;
    END
  END b1_c3
  PIN b2_c1_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 165.230 151.510 166.685 151.890 ;
        RECT 165.390 149.210 166.685 149.590 ;
        RECT 178.875 149.210 180.185 149.590 ;
        RECT 163.720 147.885 179.730 148.260 ;
        RECT 165.400 143.710 166.705 144.090 ;
        RECT 178.740 143.710 180.205 144.090 ;
        RECT 165.215 141.710 166.705 142.090 ;
      LAYER Metal2 ;
        RECT 165.520 141.000 165.875 152.085 ;
        RECT 179.030 143.430 179.360 149.625 ;
    END
  END b2_c1_not
  PIN b2_c1
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 188.925 151.610 190.205 151.990 ;
        RECT 175.425 149.210 176.610 149.590 ;
        RECT 188.925 149.210 189.940 149.590 ;
        RECT 163.720 146.530 189.950 146.920 ;
        RECT 175.405 143.710 176.765 144.090 ;
        RECT 188.905 143.710 190.085 144.090 ;
        RECT 188.905 141.710 189.980 142.090 ;
      LAYER Metal2 ;
        RECT 176.045 149.575 176.355 149.605 ;
        RECT 176.045 143.475 176.360 149.575 ;
        RECT 189.545 141.480 189.875 152.175 ;
    END
  END b2_c1
  PIN b2_c2_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 165.290 131.705 166.745 132.085 ;
        RECT 165.450 129.405 166.745 129.785 ;
        RECT 178.935 129.405 180.245 129.785 ;
        RECT 163.780 128.080 179.790 128.455 ;
        RECT 165.460 123.905 166.765 124.285 ;
        RECT 178.800 123.905 180.265 124.285 ;
        RECT 165.275 121.905 166.765 122.285 ;
      LAYER Metal2 ;
        RECT 165.580 121.195 165.935 132.280 ;
        RECT 179.090 123.625 179.420 129.820 ;
    END
  END b2_c2_not
  PIN b2_c2
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 188.985 131.805 190.265 132.185 ;
        RECT 175.485 129.405 176.670 129.785 ;
        RECT 188.985 129.405 190.000 129.785 ;
        RECT 163.780 126.725 190.010 127.115 ;
        RECT 175.465 123.905 176.825 124.285 ;
        RECT 188.965 123.905 190.145 124.285 ;
        RECT 188.965 121.905 190.040 122.285 ;
      LAYER Metal2 ;
        RECT 176.105 129.770 176.415 129.800 ;
        RECT 176.105 123.670 176.420 129.770 ;
        RECT 189.605 121.675 189.935 132.370 ;
    END
  END b2_c2
  PIN b2_c3_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 165.220 111.935 166.675 112.315 ;
        RECT 165.380 109.635 166.675 110.015 ;
        RECT 178.865 109.635 180.175 110.015 ;
        RECT 163.710 108.310 179.720 108.685 ;
        RECT 165.390 104.135 166.695 104.515 ;
        RECT 178.730 104.135 180.195 104.515 ;
        RECT 165.205 102.135 166.695 102.515 ;
      LAYER Metal2 ;
        RECT 165.510 101.425 165.865 112.510 ;
        RECT 179.020 103.855 179.350 110.050 ;
    END
  END b2_c3_not
  PIN b2_c3
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 188.915 112.035 190.195 112.415 ;
        RECT 175.415 109.635 176.600 110.015 ;
        RECT 188.915 109.635 189.930 110.015 ;
        RECT 163.710 106.955 189.940 107.345 ;
        RECT 175.395 104.135 176.755 104.515 ;
        RECT 188.895 104.135 190.075 104.515 ;
        RECT 188.895 102.135 189.970 102.515 ;
      LAYER Metal2 ;
        RECT 176.035 110.000 176.345 110.030 ;
        RECT 176.035 103.900 176.350 110.000 ;
        RECT 189.535 101.905 189.865 112.600 ;
    END
  END b2_c3
  PIN b2_c4_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 165.250 92.210 166.705 92.590 ;
        RECT 165.410 89.910 166.705 90.290 ;
        RECT 178.895 89.910 180.205 90.290 ;
        RECT 163.740 88.585 179.750 88.960 ;
        RECT 165.420 84.410 166.725 84.790 ;
        RECT 178.760 84.410 180.225 84.790 ;
        RECT 165.235 82.410 166.725 82.790 ;
      LAYER Metal2 ;
        RECT 165.540 81.700 165.895 92.785 ;
        RECT 179.050 84.130 179.380 90.325 ;
    END
  END b2_c4_not
  PIN b0_c5_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -30.920 92.200 -29.465 92.580 ;
        RECT -30.760 89.900 -29.465 90.280 ;
        RECT -17.275 89.900 -15.965 90.280 ;
        RECT -32.430 88.575 -16.420 88.950 ;
        RECT -30.750 84.400 -29.445 84.780 ;
        RECT -17.410 84.400 -15.945 84.780 ;
        RECT -30.935 82.400 -29.445 82.780 ;
      LAYER Metal2 ;
        RECT -30.630 81.690 -30.275 92.775 ;
        RECT -17.120 84.120 -16.790 90.315 ;
    END
  END b0_c5_not
  PIN b0_c5
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -7.225 92.300 -5.945 92.680 ;
        RECT -20.725 89.900 -19.540 90.280 ;
        RECT -7.225 89.900 -6.210 90.280 ;
        RECT -32.430 87.220 -6.200 87.610 ;
        RECT -20.745 84.400 -19.385 84.780 ;
        RECT -7.245 84.400 -6.065 84.780 ;
        RECT -7.245 82.400 -6.170 82.780 ;
      LAYER Metal2 ;
        RECT -20.105 90.265 -19.795 90.295 ;
        RECT -20.105 84.165 -19.790 90.265 ;
        RECT -6.605 82.170 -6.275 92.865 ;
    END
  END b0_c5
  PIN b0_c6_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -30.990 72.370 -29.535 72.750 ;
        RECT -30.830 70.070 -29.535 70.450 ;
        RECT -17.345 70.070 -16.035 70.450 ;
        RECT -32.500 68.745 -16.490 69.120 ;
        RECT -30.820 64.570 -29.515 64.950 ;
        RECT -17.480 64.570 -16.015 64.950 ;
        RECT -31.005 62.570 -29.515 62.950 ;
      LAYER Metal2 ;
        RECT -30.700 61.860 -30.345 72.945 ;
        RECT -17.190 64.290 -16.860 70.485 ;
    END
  END b0_c6_not
  PIN b0_c6
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -7.295 72.470 -6.015 72.850 ;
        RECT -20.795 70.070 -19.610 70.450 ;
        RECT -7.295 70.070 -6.280 70.450 ;
        RECT -32.500 67.390 -6.270 67.780 ;
        RECT -20.815 64.570 -19.455 64.950 ;
        RECT -7.315 64.570 -6.135 64.950 ;
        RECT -7.315 62.570 -6.240 62.950 ;
      LAYER Metal2 ;
        RECT -20.175 70.435 -19.865 70.465 ;
        RECT -20.175 64.335 -19.860 70.435 ;
        RECT -6.675 62.340 -6.345 73.035 ;
    END
  END b0_c6
  PIN b0_c7_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -30.920 52.650 -29.465 53.030 ;
        RECT -30.760 50.350 -29.465 50.730 ;
        RECT -17.275 50.350 -15.965 50.730 ;
        RECT -32.430 49.025 -16.420 49.400 ;
        RECT -30.750 44.850 -29.445 45.230 ;
        RECT -17.410 44.850 -15.945 45.230 ;
        RECT -30.935 42.850 -29.445 43.230 ;
      LAYER Metal2 ;
        RECT -30.630 42.140 -30.275 53.225 ;
        RECT -17.120 44.570 -16.790 50.765 ;
    END
  END b0_c7_not
  PIN b0_c7
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -7.225 52.750 -5.945 53.130 ;
        RECT -20.725 50.350 -19.540 50.730 ;
        RECT -7.225 50.350 -6.210 50.730 ;
        RECT -32.430 47.670 -6.200 48.060 ;
        RECT -20.745 44.850 -19.385 45.230 ;
        RECT -7.245 44.850 -6.065 45.230 ;
        RECT -7.245 42.850 -6.170 43.230 ;
      LAYER Metal2 ;
        RECT -20.105 50.715 -19.795 50.745 ;
        RECT -20.105 44.615 -19.790 50.715 ;
        RECT -6.605 42.620 -6.275 53.315 ;
    END
  END b0_c7
  PIN b2_c4
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 188.945 92.310 190.225 92.690 ;
        RECT 175.445 89.910 176.630 90.290 ;
        RECT 188.945 89.910 189.960 90.290 ;
        RECT 163.740 87.230 189.970 87.620 ;
        RECT 175.425 84.410 176.785 84.790 ;
        RECT 188.925 84.410 190.105 84.790 ;
        RECT 188.925 82.410 190.000 82.790 ;
      LAYER Metal2 ;
        RECT 176.065 90.275 176.375 90.305 ;
        RECT 176.065 84.175 176.380 90.275 ;
        RECT 189.565 82.180 189.895 92.875 ;
    END
  END b2_c4
  PIN b2_c5_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 165.180 72.380 166.635 72.760 ;
        RECT 165.340 70.080 166.635 70.460 ;
        RECT 178.825 70.080 180.135 70.460 ;
        RECT 163.670 68.755 179.680 69.130 ;
        RECT 165.350 64.580 166.655 64.960 ;
        RECT 178.690 64.580 180.155 64.960 ;
        RECT 165.165 62.580 166.655 62.960 ;
      LAYER Metal2 ;
        RECT 165.470 61.870 165.825 72.955 ;
        RECT 178.980 64.300 179.310 70.495 ;
    END
  END b2_c5_not
  PIN b2_c5
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 188.875 72.480 190.155 72.860 ;
        RECT 175.375 70.080 176.560 70.460 ;
        RECT 188.875 70.080 189.890 70.460 ;
        RECT 163.670 67.400 189.900 67.790 ;
        RECT 175.355 64.580 176.715 64.960 ;
        RECT 188.855 64.580 190.035 64.960 ;
        RECT 188.855 62.580 189.930 62.960 ;
      LAYER Metal2 ;
        RECT 175.995 70.445 176.305 70.475 ;
        RECT 175.995 64.345 176.310 70.445 ;
        RECT 189.495 62.350 189.825 73.045 ;
    END
  END b2_c5
  PIN b2_c6_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 165.250 52.660 166.705 53.040 ;
        RECT 165.410 50.360 166.705 50.740 ;
        RECT 178.895 50.360 180.205 50.740 ;
        RECT 163.740 49.035 179.750 49.410 ;
        RECT 165.420 44.860 166.725 45.240 ;
        RECT 178.760 44.860 180.225 45.240 ;
        RECT 165.235 42.860 166.725 43.240 ;
      LAYER Metal2 ;
        RECT 165.540 42.150 165.895 53.235 ;
        RECT 179.050 44.580 179.380 50.775 ;
    END
  END b2_c6_not
  PIN b2_c6
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 188.945 52.760 190.225 53.140 ;
        RECT 175.445 50.360 176.630 50.740 ;
        RECT 188.945 50.360 189.960 50.740 ;
        RECT 163.740 47.680 189.970 48.070 ;
        RECT 175.425 44.860 176.785 45.240 ;
        RECT 188.925 44.860 190.105 45.240 ;
        RECT 188.925 42.860 190.000 43.240 ;
      LAYER Metal2 ;
        RECT 176.065 50.725 176.375 50.755 ;
        RECT 176.065 44.625 176.380 50.725 ;
        RECT 189.565 42.630 189.895 53.325 ;
    END
  END b2_c6
  PIN x0_b0_f
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 81.980 10.895 82.360 11.275 ;
        RECT 80.380 10.380 81.580 10.670 ;
        RECT 72.645 8.210 81.575 8.510 ;
        RECT 81.170 4.605 82.360 4.890 ;
        RECT 80.390 3.940 80.770 4.320 ;
      LAYER Metal2 ;
        RECT 80.430 3.930 80.730 10.740 ;
        RECT 81.220 4.525 81.530 10.715 ;
        RECT 82.015 4.455 82.315 11.285 ;
    END
  END x0_b0_f
  PIN b2_c7_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 165.225 32.930 166.680 33.310 ;
        RECT 165.385 30.630 166.680 31.010 ;
        RECT 178.870 30.630 180.180 31.010 ;
        RECT 163.715 29.305 179.725 29.680 ;
        RECT 165.395 25.130 166.700 25.510 ;
        RECT 178.735 25.130 180.200 25.510 ;
        RECT 165.210 23.130 166.700 23.510 ;
      LAYER Metal2 ;
        RECT 165.515 22.420 165.870 33.505 ;
        RECT 179.025 24.850 179.355 31.045 ;
    END
  END b2_c7_not
  PIN b2_c7
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 188.920 33.030 190.200 33.410 ;
        RECT 175.420 30.630 176.605 31.010 ;
        RECT 188.920 30.630 189.935 31.010 ;
        RECT 163.715 27.950 189.945 28.340 ;
        RECT 175.400 25.130 176.760 25.510 ;
        RECT 188.900 25.130 190.080 25.510 ;
        RECT 188.900 23.130 189.975 23.510 ;
      LAYER Metal2 ;
        RECT 176.040 30.995 176.350 31.025 ;
        RECT 176.040 24.895 176.355 30.995 ;
        RECT 189.540 22.900 189.870 33.595 ;
    END
  END b2_c7
  PIN b1_c4_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -81.245 92.120 -79.790 92.500 ;
        RECT -81.085 89.820 -79.790 90.200 ;
        RECT -67.600 89.820 -66.290 90.200 ;
        RECT -82.755 88.495 -66.745 88.870 ;
        RECT -81.075 84.320 -79.770 84.700 ;
        RECT -67.735 84.320 -66.270 84.700 ;
        RECT -81.260 82.320 -79.770 82.700 ;
      LAYER Metal2 ;
        RECT -80.955 81.610 -80.600 92.695 ;
        RECT -67.445 84.040 -67.115 90.235 ;
    END
  END b1_c4_not
  PIN b1_c4
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -57.550 92.220 -56.270 92.600 ;
        RECT -71.050 89.820 -69.865 90.200 ;
        RECT -57.550 89.820 -56.535 90.200 ;
        RECT -82.755 87.140 -56.525 87.530 ;
        RECT -71.070 84.320 -69.710 84.700 ;
        RECT -57.570 84.320 -56.390 84.700 ;
        RECT -57.570 82.320 -56.495 82.700 ;
      LAYER Metal2 ;
        RECT -70.430 90.185 -70.120 90.215 ;
        RECT -70.430 84.085 -70.115 90.185 ;
        RECT -56.930 82.090 -56.600 92.785 ;
    END
  END b1_c4
  PIN b1_c5_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -81.315 72.290 -79.860 72.670 ;
        RECT -81.155 69.990 -79.860 70.370 ;
        RECT -67.670 69.990 -66.360 70.370 ;
        RECT -82.825 68.665 -66.815 69.040 ;
        RECT -81.145 64.490 -79.840 64.870 ;
        RECT -67.805 64.490 -66.340 64.870 ;
        RECT -81.330 62.490 -79.840 62.870 ;
      LAYER Metal2 ;
        RECT -81.025 61.780 -80.670 72.865 ;
        RECT -67.515 64.210 -67.185 70.405 ;
    END
  END b1_c5_not
  PIN b1_c5
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -57.620 72.390 -56.340 72.770 ;
        RECT -71.120 69.990 -69.935 70.370 ;
        RECT -57.620 69.990 -56.605 70.370 ;
        RECT -82.825 67.310 -56.595 67.700 ;
        RECT -71.140 64.490 -69.780 64.870 ;
        RECT -57.640 64.490 -56.460 64.870 ;
        RECT -57.640 62.490 -56.565 62.870 ;
      LAYER Metal2 ;
        RECT -70.500 70.355 -70.190 70.385 ;
        RECT -70.500 64.255 -70.185 70.355 ;
        RECT -57.000 62.260 -56.670 72.955 ;
    END
  END b1_c5
  PIN b1_c6_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -81.245 52.570 -79.790 52.950 ;
        RECT -81.085 50.270 -79.790 50.650 ;
        RECT -67.600 50.270 -66.290 50.650 ;
        RECT -82.755 48.945 -66.745 49.320 ;
        RECT -81.075 44.770 -79.770 45.150 ;
        RECT -67.735 44.770 -66.270 45.150 ;
        RECT -81.260 42.770 -79.770 43.150 ;
      LAYER Metal2 ;
        RECT -80.955 42.060 -80.600 53.145 ;
        RECT -67.445 44.490 -67.115 50.685 ;
    END
  END b1_c6_not
  PIN b1_c6
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -57.550 52.670 -56.270 53.050 ;
        RECT -71.050 50.270 -69.865 50.650 ;
        RECT -57.550 50.270 -56.535 50.650 ;
        RECT -82.755 47.590 -56.525 47.980 ;
        RECT -71.070 44.770 -69.710 45.150 ;
        RECT -57.570 44.770 -56.390 45.150 ;
        RECT -57.570 42.770 -56.495 43.150 ;
      LAYER Metal2 ;
        RECT -70.430 50.635 -70.120 50.665 ;
        RECT -70.430 44.535 -70.115 50.635 ;
        RECT -56.930 42.540 -56.600 53.235 ;
    END
  END b1_c6
  PIN b1_c7_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -81.240 32.760 -79.785 33.140 ;
        RECT -81.080 30.460 -79.785 30.840 ;
        RECT -67.595 30.460 -66.285 30.840 ;
        RECT -82.750 29.135 -66.740 29.510 ;
        RECT -81.070 24.960 -79.765 25.340 ;
        RECT -67.730 24.960 -66.265 25.340 ;
        RECT -81.255 22.960 -79.765 23.340 ;
      LAYER Metal2 ;
        RECT -80.950 22.250 -80.595 33.335 ;
        RECT -67.440 24.680 -67.110 30.875 ;
    END
  END b1_c7_not
  PIN b1_c7
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT -57.545 32.860 -56.265 33.240 ;
        RECT -71.045 30.460 -69.860 30.840 ;
        RECT -57.545 30.460 -56.530 30.840 ;
        RECT -82.750 27.780 -56.520 28.170 ;
        RECT -71.065 24.960 -69.705 25.340 ;
        RECT -57.565 24.960 -56.385 25.340 ;
        RECT -57.565 22.960 -56.490 23.340 ;
      LAYER Metal2 ;
        RECT -70.425 30.825 -70.115 30.855 ;
        RECT -70.425 24.725 -70.110 30.825 ;
        RECT -56.925 22.730 -56.595 33.425 ;
    END
  END b1_c7
  PIN x0_b0_f_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 75.520 11.115 78.930 11.495 ;
        RECT 87.300 10.445 87.680 10.825 ;
        RECT 72.615 7.675 78.955 7.945 ;
        RECT 78.530 6.415 84.920 6.705 ;
        RECT 75.510 4.500 75.890 4.880 ;
        RECT 84.510 3.775 87.690 4.095 ;
      LAYER Metal2 ;
        RECT 75.555 4.445 75.855 11.485 ;
        RECT 78.580 6.315 78.905 11.475 ;
        RECT 84.590 3.715 84.870 6.750 ;
        RECT 87.340 3.670 87.640 10.825 ;
    END
  END x0_b0_f_not
  PIN b4_c5
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 581.585 72.485 582.865 72.865 ;
        RECT 568.085 70.085 569.270 70.465 ;
        RECT 581.585 70.085 582.600 70.465 ;
        RECT 556.380 67.405 582.610 67.795 ;
        RECT 568.065 64.585 569.425 64.965 ;
        RECT 581.565 64.585 582.745 64.965 ;
        RECT 581.565 62.585 582.640 62.965 ;
      LAYER Metal2 ;
        RECT 568.705 70.450 569.015 70.480 ;
        RECT 568.705 64.350 569.020 70.450 ;
        RECT 582.205 62.355 582.535 73.050 ;
    END
  END b4_c5
  PIN b3_c7
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 385.310 32.990 386.590 33.370 ;
        RECT 371.810 30.590 372.995 30.970 ;
        RECT 385.310 30.590 386.325 30.970 ;
        RECT 360.105 27.910 386.335 28.300 ;
        RECT 371.790 25.090 373.150 25.470 ;
        RECT 385.290 25.090 386.470 25.470 ;
        RECT 385.290 23.090 386.365 23.470 ;
      LAYER Metal2 ;
        RECT 372.430 30.955 372.740 30.985 ;
        RECT 372.430 24.855 372.745 30.955 ;
        RECT 385.930 22.860 386.260 33.555 ;
    END
  END b3_c7
  PIN b4_c7_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 557.935 32.935 559.390 33.315 ;
        RECT 558.095 30.635 559.390 31.015 ;
        RECT 571.580 30.635 572.890 31.015 ;
        RECT 556.425 29.310 572.435 29.685 ;
        RECT 558.105 25.135 559.410 25.515 ;
        RECT 571.445 25.135 572.910 25.515 ;
        RECT 557.920 23.135 559.410 23.515 ;
      LAYER Metal2 ;
        RECT 558.225 22.425 558.580 33.510 ;
        RECT 571.735 24.855 572.065 31.050 ;
    END
  END b4_c7_not
  PIN b4_c7
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 581.630 33.035 582.910 33.415 ;
        RECT 568.130 30.635 569.315 31.015 ;
        RECT 581.630 30.635 582.645 31.015 ;
        RECT 556.425 27.955 582.655 28.345 ;
        RECT 568.110 25.135 569.470 25.515 ;
        RECT 581.610 25.135 582.790 25.515 ;
        RECT 581.610 23.135 582.685 23.515 ;
      LAYER Metal2 ;
        RECT 568.750 31.000 569.060 31.030 ;
        RECT 568.750 24.900 569.065 31.000 ;
        RECT 582.250 22.905 582.580 33.600 ;
    END
  END b4_c7
  PIN b3_c4_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 361.640 92.170 363.095 92.550 ;
        RECT 361.800 89.870 363.095 90.250 ;
        RECT 375.285 89.870 376.595 90.250 ;
        RECT 360.130 88.545 376.140 88.920 ;
        RECT 361.810 84.370 363.115 84.750 ;
        RECT 375.150 84.370 376.615 84.750 ;
        RECT 361.625 82.370 363.115 82.750 ;
      LAYER Metal2 ;
        RECT 361.930 81.660 362.285 92.745 ;
        RECT 375.440 84.090 375.770 90.285 ;
    END
  END b3_c4_not
  PIN b3_c4
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 385.335 92.270 386.615 92.650 ;
        RECT 371.835 89.870 373.020 90.250 ;
        RECT 385.335 89.870 386.350 90.250 ;
        RECT 360.130 87.190 386.360 87.580 ;
        RECT 371.815 84.370 373.175 84.750 ;
        RECT 385.315 84.370 386.495 84.750 ;
        RECT 385.315 82.370 386.390 82.750 ;
      LAYER Metal2 ;
        RECT 372.455 90.235 372.765 90.265 ;
        RECT 372.455 84.135 372.770 90.235 ;
        RECT 385.955 82.140 386.285 92.835 ;
    END
  END b3_c4
  PIN b3_c5_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 361.570 72.340 363.025 72.720 ;
        RECT 361.730 70.040 363.025 70.420 ;
        RECT 375.215 70.040 376.525 70.420 ;
        RECT 360.060 68.715 376.070 69.090 ;
        RECT 361.740 64.540 363.045 64.920 ;
        RECT 375.080 64.540 376.545 64.920 ;
        RECT 361.555 62.540 363.045 62.920 ;
      LAYER Metal2 ;
        RECT 361.860 61.830 362.215 72.915 ;
        RECT 375.370 64.260 375.700 70.455 ;
    END
  END b3_c5_not
  PIN b3_c5
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 385.265 72.440 386.545 72.820 ;
        RECT 371.765 70.040 372.950 70.420 ;
        RECT 385.265 70.040 386.280 70.420 ;
        RECT 360.060 67.360 386.290 67.750 ;
        RECT 371.745 64.540 373.105 64.920 ;
        RECT 385.245 64.540 386.425 64.920 ;
        RECT 385.245 62.540 386.320 62.920 ;
      LAYER Metal2 ;
        RECT 372.385 70.405 372.695 70.435 ;
        RECT 372.385 64.305 372.700 70.405 ;
        RECT 385.885 62.310 386.215 73.005 ;
    END
  END b3_c5
  PIN b3_c6_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 361.640 52.620 363.095 53.000 ;
        RECT 361.800 50.320 363.095 50.700 ;
        RECT 375.285 50.320 376.595 50.700 ;
        RECT 360.130 48.995 376.140 49.370 ;
        RECT 361.810 44.820 363.115 45.200 ;
        RECT 375.150 44.820 376.615 45.200 ;
        RECT 361.625 42.820 363.115 43.200 ;
      LAYER Metal2 ;
        RECT 361.930 42.110 362.285 53.195 ;
        RECT 375.440 44.540 375.770 50.735 ;
    END
  END b3_c6_not
  PIN x1_b0_f
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 278.345 10.895 278.725 11.275 ;
        RECT 276.745 10.380 277.945 10.670 ;
        RECT 269.010 8.210 277.940 8.510 ;
        RECT 277.535 4.605 278.725 4.890 ;
        RECT 276.755 3.940 277.135 4.320 ;
      LAYER Metal2 ;
        RECT 276.795 3.930 277.095 10.740 ;
        RECT 277.585 4.525 277.895 10.715 ;
        RECT 278.380 4.455 278.680 11.285 ;
    END
  END x1_b0_f
  PIN x1_b0_f_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 271.885 11.115 275.295 11.495 ;
        RECT 283.665 10.445 284.045 10.825 ;
        RECT 268.980 7.675 275.320 7.945 ;
        RECT 274.895 6.415 281.285 6.705 ;
        RECT 271.875 4.500 272.255 4.880 ;
        RECT 280.875 3.775 284.055 4.095 ;
      LAYER Metal2 ;
        RECT 271.920 4.445 272.220 11.485 ;
        RECT 274.945 6.315 275.270 11.475 ;
        RECT 280.955 3.715 281.235 6.750 ;
        RECT 283.705 3.670 284.005 10.825 ;
    END
  END x1_b0_f_not
  PIN x2_b0_f
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 474.745 10.845 475.125 11.225 ;
        RECT 473.145 10.330 474.345 10.620 ;
        RECT 465.410 8.160 474.340 8.460 ;
        RECT 473.935 4.555 475.125 4.840 ;
        RECT 473.155 3.890 473.535 4.270 ;
      LAYER Metal2 ;
        RECT 473.195 3.880 473.495 10.690 ;
        RECT 473.985 4.475 474.295 10.665 ;
        RECT 474.780 4.405 475.080 11.235 ;
    END
  END x2_b0_f
  PIN x2_b0_f_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 468.285 11.065 471.695 11.445 ;
        RECT 480.065 10.395 480.445 10.775 ;
        RECT 465.380 7.625 471.720 7.895 ;
        RECT 471.295 6.365 477.685 6.655 ;
        RECT 468.275 4.450 468.655 4.830 ;
        RECT 477.275 3.725 480.455 4.045 ;
      LAYER Metal2 ;
        RECT 468.320 4.395 468.620 11.435 ;
        RECT 471.345 6.265 471.670 11.425 ;
        RECT 477.355 3.665 477.635 6.700 ;
        RECT 480.105 3.620 480.405 10.775 ;
    END
  END x2_b0_f_not
  PIN b4_c6_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 557.960 52.665 559.415 53.045 ;
        RECT 558.120 50.365 559.415 50.745 ;
        RECT 571.605 50.365 572.915 50.745 ;
        RECT 556.450 49.040 572.460 49.415 ;
        RECT 558.130 44.865 559.435 45.245 ;
        RECT 571.470 44.865 572.935 45.245 ;
        RECT 557.945 42.865 559.435 43.245 ;
      LAYER Metal2 ;
        RECT 558.250 42.155 558.605 53.240 ;
        RECT 571.760 44.585 572.090 50.780 ;
    END
  END b4_c6_not
  PIN b4_c6
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 581.655 52.765 582.935 53.145 ;
        RECT 568.155 50.365 569.340 50.745 ;
        RECT 581.655 50.365 582.670 50.745 ;
        RECT 556.450 47.685 582.680 48.075 ;
        RECT 568.135 44.865 569.495 45.245 ;
        RECT 581.635 44.865 582.815 45.245 ;
        RECT 581.635 42.865 582.710 43.245 ;
      LAYER Metal2 ;
        RECT 568.775 50.730 569.085 50.760 ;
        RECT 568.775 44.630 569.090 50.730 ;
        RECT 582.275 42.635 582.605 53.330 ;
    END
  END b4_c6
  PIN b3_c6
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 385.335 52.720 386.615 53.100 ;
        RECT 371.835 50.320 373.020 50.700 ;
        RECT 385.335 50.320 386.350 50.700 ;
        RECT 360.130 47.640 386.360 48.030 ;
        RECT 371.815 44.820 373.175 45.200 ;
        RECT 385.315 44.820 386.495 45.200 ;
        RECT 385.315 42.820 386.390 43.200 ;
      LAYER Metal2 ;
        RECT 372.455 50.685 372.765 50.715 ;
        RECT 372.455 44.585 372.770 50.685 ;
        RECT 385.955 42.590 386.285 53.285 ;
    END
  END b3_c6
  PIN b3_c7_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 361.615 32.890 363.070 33.270 ;
        RECT 361.775 30.590 363.070 30.970 ;
        RECT 375.260 30.590 376.570 30.970 ;
        RECT 360.105 29.265 376.115 29.640 ;
        RECT 361.785 25.090 363.090 25.470 ;
        RECT 375.125 25.090 376.590 25.470 ;
        RECT 361.600 23.090 363.090 23.470 ;
      LAYER Metal2 ;
        RECT 361.905 22.380 362.260 33.465 ;
        RECT 375.415 24.810 375.745 31.005 ;
    END
  END b3_c7_not
  PIN b4_c4_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 557.960 92.215 559.415 92.595 ;
        RECT 558.120 89.915 559.415 90.295 ;
        RECT 571.605 89.915 572.915 90.295 ;
        RECT 556.450 88.590 572.460 88.965 ;
        RECT 558.130 84.415 559.435 84.795 ;
        RECT 571.470 84.415 572.935 84.795 ;
        RECT 557.945 82.415 559.435 82.795 ;
      LAYER Metal2 ;
        RECT 558.250 81.705 558.605 92.790 ;
        RECT 571.760 84.135 572.090 90.330 ;
    END
  END b4_c4_not
  PIN b4_c4
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 581.655 92.315 582.935 92.695 ;
        RECT 568.155 89.915 569.340 90.295 ;
        RECT 581.655 89.915 582.670 90.295 ;
        RECT 556.450 87.235 582.680 87.625 ;
        RECT 568.135 84.415 569.495 84.795 ;
        RECT 581.635 84.415 582.815 84.795 ;
        RECT 581.635 82.415 582.710 82.795 ;
      LAYER Metal2 ;
        RECT 568.775 90.280 569.085 90.310 ;
        RECT 568.775 84.180 569.090 90.280 ;
        RECT 582.275 82.185 582.605 92.880 ;
    END
  END b4_c4
  PIN b4_c5_not
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 557.890 72.385 559.345 72.765 ;
        RECT 558.050 70.085 559.345 70.465 ;
        RECT 571.535 70.085 572.845 70.465 ;
        RECT 556.380 68.760 572.390 69.135 ;
        RECT 558.060 64.585 559.365 64.965 ;
        RECT 571.400 64.585 572.865 64.965 ;
        RECT 557.875 62.585 559.365 62.965 ;
      LAYER Metal2 ;
        RECT 558.180 61.875 558.535 72.960 ;
        RECT 571.690 64.305 572.020 70.500 ;
    END
  END b4_c5_not
  PIN p15_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 1264.325 10.830 1264.705 11.210 ;
        RECT 1261.250 10.360 1263.840 10.710 ;
        RECT 1263.435 7.895 1266.510 8.170 ;
        RECT 1263.450 4.470 1264.760 4.790 ;
        RECT 1261.260 3.915 1261.640 4.295 ;
      LAYER Metal2 ;
        RECT 1261.300 3.825 1261.600 10.765 ;
        RECT 1263.510 4.400 1263.815 10.760 ;
        RECT 1264.360 4.400 1264.660 11.220 ;
        RECT 1266.090 7.840 1266.470 8.220 ;
      LAYER Metal3 ;
        RECT 1266.055 7.885 1269.460 8.170 ;
    END
  END p15_not
  PIN b4_r0_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 667.720 171.120 668.920 171.500 ;
        RECT 667.720 168.820 670.980 169.200 ;
        RECT 668.385 166.905 690.940 167.245 ;
        RECT 692.050 166.915 706.695 167.215 ;
        RECT 667.700 163.320 671.000 163.700 ;
        RECT 695.075 163.240 697.995 163.540 ;
        RECT 701.540 163.225 704.910 163.525 ;
        RECT 667.700 161.320 668.985 161.700 ;
      LAYER Metal2 ;
        RECT 668.545 160.590 668.860 171.640 ;
        RECT 690.520 166.835 690.940 167.295 ;
        RECT 692.020 166.830 692.440 167.290 ;
        RECT 695.110 163.190 695.410 167.250 ;
        RECT 701.600 163.175 701.880 167.265 ;
        RECT 706.365 166.785 706.670 172.260 ;
      LAYER Metal3 ;
        RECT 706.320 171.750 721.800 172.205 ;
        RECT 690.490 166.885 692.515 167.270 ;
    END
  END b4_r0_b_not
  PIN b4_r1_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 667.520 151.395 668.720 151.775 ;
        RECT 667.520 149.095 670.780 149.475 ;
        RECT 668.185 147.180 690.740 147.520 ;
        RECT 691.850 147.190 706.495 147.490 ;
        RECT 667.500 143.595 670.800 143.975 ;
        RECT 694.875 143.515 697.795 143.815 ;
        RECT 701.340 143.500 704.710 143.800 ;
        RECT 667.500 141.595 668.785 141.975 ;
      LAYER Metal2 ;
        RECT 668.345 140.865 668.660 151.915 ;
        RECT 690.320 147.110 690.740 147.570 ;
        RECT 691.820 147.105 692.240 147.565 ;
        RECT 694.910 143.465 695.210 147.525 ;
        RECT 701.400 143.450 701.680 147.540 ;
        RECT 706.165 147.060 706.470 152.535 ;
      LAYER Metal3 ;
        RECT 706.120 152.025 721.600 152.480 ;
        RECT 690.290 147.160 692.315 147.545 ;
    END
  END b4_r1_b_not
  PIN b4_r0_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 687.245 171.220 688.480 171.600 ;
        RECT 685.220 168.820 688.480 169.200 ;
        RECT 692.650 167.660 706.265 167.960 ;
        RECT 693.845 165.005 697.975 165.305 ;
        RECT 700.350 164.955 704.850 165.265 ;
        RECT 687.105 163.960 691.050 164.295 ;
        RECT 685.200 163.320 688.500 163.700 ;
        RECT 687.015 161.320 688.500 161.700 ;
      LAYER Metal2 ;
        RECT 687.330 161.075 687.645 171.760 ;
        RECT 690.655 163.945 691.035 164.325 ;
        RECT 692.720 163.920 693.030 168.040 ;
        RECT 705.790 167.615 706.085 172.985 ;
      LAYER Metal3 ;
        RECT 705.790 172.530 721.810 172.940 ;
        RECT 690.655 163.935 693.135 164.335 ;
    END
  END b4_r0_b
  PIN b4_r1_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 687.045 151.495 688.280 151.875 ;
        RECT 685.020 149.095 688.280 149.475 ;
        RECT 692.450 147.935 706.065 148.235 ;
        RECT 693.645 145.280 697.775 145.580 ;
        RECT 700.150 145.230 704.650 145.540 ;
        RECT 686.905 144.235 690.850 144.570 ;
        RECT 685.000 143.595 688.300 143.975 ;
        RECT 686.815 141.595 688.300 141.975 ;
      LAYER Metal2 ;
        RECT 687.130 141.350 687.445 152.035 ;
        RECT 690.455 144.220 690.835 144.600 ;
        RECT 692.520 144.195 692.830 148.315 ;
        RECT 705.590 147.890 705.885 153.260 ;
      LAYER Metal3 ;
        RECT 705.590 152.805 721.610 153.215 ;
        RECT 690.455 144.210 692.935 144.610 ;
    END
  END b4_r1_b
  PIN b4_r2_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 667.675 131.750 668.875 132.130 ;
        RECT 667.675 129.450 670.935 129.830 ;
        RECT 668.340 127.535 690.895 127.875 ;
        RECT 692.005 127.545 706.650 127.845 ;
        RECT 667.655 123.950 670.955 124.330 ;
        RECT 695.030 123.870 697.950 124.170 ;
        RECT 701.495 123.855 704.865 124.155 ;
        RECT 667.655 121.950 668.940 122.330 ;
      LAYER Metal2 ;
        RECT 668.500 121.220 668.815 132.270 ;
        RECT 690.475 127.465 690.895 127.925 ;
        RECT 691.975 127.460 692.395 127.920 ;
        RECT 695.065 123.820 695.365 127.880 ;
        RECT 701.555 123.805 701.835 127.895 ;
        RECT 706.320 127.415 706.625 132.890 ;
      LAYER Metal3 ;
        RECT 706.275 132.380 721.755 132.835 ;
        RECT 690.445 127.515 692.470 127.900 ;
    END
  END b4_r2_b_not
  PIN b4_r2_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 687.200 131.850 688.435 132.230 ;
        RECT 685.175 129.450 688.435 129.830 ;
        RECT 692.605 128.290 706.220 128.590 ;
        RECT 693.800 125.635 697.930 125.935 ;
        RECT 700.305 125.585 704.805 125.895 ;
        RECT 687.060 124.590 691.005 124.925 ;
        RECT 685.155 123.950 688.455 124.330 ;
        RECT 686.970 121.950 688.455 122.330 ;
      LAYER Metal2 ;
        RECT 687.285 121.705 687.600 132.390 ;
        RECT 690.610 124.575 690.990 124.955 ;
        RECT 692.675 124.550 692.985 128.670 ;
        RECT 705.745 128.245 706.040 133.615 ;
      LAYER Metal3 ;
        RECT 705.745 133.160 721.765 133.570 ;
        RECT 690.610 124.565 693.090 124.965 ;
    END
  END b4_r2_b
  PIN b4_r3_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 667.675 111.955 668.875 112.335 ;
        RECT 667.675 109.655 670.935 110.035 ;
        RECT 668.340 107.740 690.895 108.080 ;
        RECT 692.005 107.750 706.650 108.050 ;
        RECT 667.655 104.155 670.955 104.535 ;
        RECT 695.030 104.075 697.950 104.375 ;
        RECT 701.495 104.060 704.865 104.360 ;
        RECT 667.655 102.155 668.940 102.535 ;
      LAYER Metal2 ;
        RECT 668.500 101.425 668.815 112.475 ;
        RECT 690.475 107.670 690.895 108.130 ;
        RECT 691.975 107.665 692.395 108.125 ;
        RECT 695.065 104.025 695.365 108.085 ;
        RECT 701.555 104.010 701.835 108.100 ;
        RECT 706.320 107.620 706.625 113.095 ;
      LAYER Metal3 ;
        RECT 706.275 112.585 721.755 113.040 ;
        RECT 690.445 107.720 692.470 108.105 ;
    END
  END b4_r3_b_not
  PIN b4_r3_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 687.200 112.055 688.435 112.435 ;
        RECT 685.175 109.655 688.435 110.035 ;
        RECT 692.605 108.495 706.220 108.795 ;
        RECT 693.800 105.840 697.930 106.140 ;
        RECT 700.305 105.790 704.805 106.100 ;
        RECT 687.060 104.795 691.005 105.130 ;
        RECT 685.155 104.155 688.455 104.535 ;
        RECT 686.970 102.155 688.455 102.535 ;
      LAYER Metal2 ;
        RECT 687.285 101.910 687.600 112.595 ;
        RECT 690.610 104.780 690.990 105.160 ;
        RECT 692.675 104.755 692.985 108.875 ;
        RECT 705.745 108.450 706.040 113.820 ;
      LAYER Metal3 ;
        RECT 705.745 113.365 721.765 113.775 ;
        RECT 690.610 104.770 693.090 105.170 ;
    END
  END b4_r3_b
  PIN b4_r4_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 667.595 92.200 668.795 92.580 ;
        RECT 667.595 89.900 670.855 90.280 ;
        RECT 668.260 87.985 690.815 88.325 ;
        RECT 691.925 87.995 706.570 88.295 ;
        RECT 667.575 84.400 670.875 84.780 ;
        RECT 694.950 84.320 697.870 84.620 ;
        RECT 701.415 84.305 704.785 84.605 ;
        RECT 667.575 82.400 668.860 82.780 ;
      LAYER Metal2 ;
        RECT 668.420 81.670 668.735 92.720 ;
        RECT 690.395 87.915 690.815 88.375 ;
        RECT 691.895 87.910 692.315 88.370 ;
        RECT 694.985 84.270 695.285 88.330 ;
        RECT 701.475 84.255 701.755 88.345 ;
        RECT 706.240 87.865 706.545 93.340 ;
      LAYER Metal3 ;
        RECT 706.195 92.830 721.675 93.285 ;
        RECT 690.365 87.965 692.390 88.350 ;
    END
  END b4_r4_b_not
  PIN b4_r4_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 687.120 92.300 688.355 92.680 ;
        RECT 685.095 89.900 688.355 90.280 ;
        RECT 692.525 88.740 706.140 89.040 ;
        RECT 693.720 86.085 697.850 86.385 ;
        RECT 700.225 86.035 704.725 86.345 ;
        RECT 686.980 85.040 690.925 85.375 ;
        RECT 685.075 84.400 688.375 84.780 ;
        RECT 686.890 82.400 688.375 82.780 ;
      LAYER Metal2 ;
        RECT 687.205 82.155 687.520 92.840 ;
        RECT 690.530 85.025 690.910 85.405 ;
        RECT 692.595 85.000 692.905 89.120 ;
        RECT 705.665 88.695 705.960 94.065 ;
      LAYER Metal3 ;
        RECT 705.665 93.610 721.685 94.020 ;
        RECT 690.530 85.015 693.010 85.415 ;
    END
  END b4_r4_b
  PIN b4_r5_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 667.700 72.485 668.900 72.865 ;
        RECT 667.700 70.185 670.960 70.565 ;
        RECT 668.365 68.270 690.920 68.610 ;
        RECT 692.030 68.280 706.675 68.580 ;
        RECT 667.680 64.685 670.980 65.065 ;
        RECT 695.055 64.605 697.975 64.905 ;
        RECT 701.520 64.590 704.890 64.890 ;
        RECT 667.680 62.685 668.965 63.065 ;
      LAYER Metal2 ;
        RECT 668.525 61.955 668.840 73.005 ;
        RECT 690.500 68.200 690.920 68.660 ;
        RECT 692.000 68.195 692.420 68.655 ;
        RECT 695.090 64.555 695.390 68.615 ;
        RECT 701.580 64.540 701.860 68.630 ;
        RECT 706.345 68.150 706.650 73.625 ;
      LAYER Metal3 ;
        RECT 706.300 73.115 721.780 73.570 ;
        RECT 690.470 68.250 692.495 68.635 ;
    END
  END b4_r5_b_not
  PIN b4_r5_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 687.225 72.585 688.460 72.965 ;
        RECT 685.200 70.185 688.460 70.565 ;
        RECT 692.630 69.025 706.245 69.325 ;
        RECT 693.825 66.370 697.955 66.670 ;
        RECT 700.330 66.320 704.830 66.630 ;
        RECT 687.085 65.325 691.030 65.660 ;
        RECT 685.180 64.685 688.480 65.065 ;
        RECT 686.995 62.685 688.480 63.065 ;
      LAYER Metal2 ;
        RECT 687.310 62.440 687.625 73.125 ;
        RECT 690.635 65.310 691.015 65.690 ;
        RECT 692.700 65.285 693.010 69.405 ;
        RECT 705.770 68.980 706.065 74.350 ;
      LAYER Metal3 ;
        RECT 705.770 73.895 721.790 74.305 ;
        RECT 690.635 65.300 693.115 65.700 ;
    END
  END b4_r5_b
  PIN b4_r6_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 667.700 52.515 668.900 52.895 ;
        RECT 667.700 50.215 670.960 50.595 ;
        RECT 668.365 48.300 690.920 48.640 ;
        RECT 692.030 48.310 706.675 48.610 ;
        RECT 667.680 44.715 670.980 45.095 ;
        RECT 695.055 44.635 697.975 44.935 ;
        RECT 701.520 44.620 704.890 44.920 ;
        RECT 667.680 42.715 668.965 43.095 ;
      LAYER Metal2 ;
        RECT 668.525 41.985 668.840 53.035 ;
        RECT 690.500 48.230 690.920 48.690 ;
        RECT 692.000 48.225 692.420 48.685 ;
        RECT 695.090 44.585 695.390 48.645 ;
        RECT 701.580 44.570 701.860 48.660 ;
        RECT 706.345 48.180 706.650 53.655 ;
      LAYER Metal3 ;
        RECT 706.300 53.145 721.780 53.600 ;
        RECT 690.470 48.280 692.495 48.665 ;
    END
  END b4_r6_b_not
  PIN b4_r6_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 687.225 52.615 688.460 52.995 ;
        RECT 685.200 50.215 688.460 50.595 ;
        RECT 692.630 49.055 706.245 49.355 ;
        RECT 693.825 46.400 697.955 46.700 ;
        RECT 700.330 46.350 704.830 46.660 ;
        RECT 687.085 45.355 691.030 45.690 ;
        RECT 685.180 44.715 688.480 45.095 ;
        RECT 686.995 42.715 688.480 43.095 ;
      LAYER Metal2 ;
        RECT 687.310 42.470 687.625 53.155 ;
        RECT 690.635 45.340 691.015 45.720 ;
        RECT 692.700 45.315 693.010 49.435 ;
        RECT 705.770 49.010 706.065 54.380 ;
      LAYER Metal3 ;
        RECT 705.770 53.925 721.790 54.335 ;
        RECT 690.635 45.330 693.115 45.730 ;
    END
  END b4_r6_b
  PIN b4_r7_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 667.700 32.850 668.900 33.230 ;
        RECT 667.700 30.550 670.960 30.930 ;
        RECT 668.365 28.635 690.920 28.975 ;
        RECT 692.030 28.645 706.675 28.945 ;
        RECT 667.680 25.050 670.980 25.430 ;
        RECT 695.055 24.970 697.975 25.270 ;
        RECT 701.520 24.955 704.890 25.255 ;
        RECT 667.680 23.050 668.965 23.430 ;
      LAYER Metal2 ;
        RECT 668.525 22.320 668.840 33.370 ;
        RECT 690.500 28.565 690.920 29.025 ;
        RECT 692.000 28.560 692.420 29.020 ;
        RECT 695.090 24.920 695.390 28.980 ;
        RECT 701.580 24.905 701.860 28.995 ;
        RECT 706.345 28.515 706.650 33.990 ;
      LAYER Metal3 ;
        RECT 706.300 33.480 721.780 33.935 ;
        RECT 690.470 28.615 692.495 29.000 ;
    END
  END b4_r7_b_not
  PIN b4_r7_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 687.225 32.950 688.460 33.330 ;
        RECT 685.200 30.550 688.460 30.930 ;
        RECT 692.630 29.390 706.245 29.690 ;
        RECT 693.825 26.735 697.955 27.035 ;
        RECT 700.330 26.685 704.830 26.995 ;
        RECT 687.085 25.690 691.030 26.025 ;
        RECT 685.180 25.050 688.480 25.430 ;
        RECT 686.995 23.050 688.480 23.430 ;
      LAYER Metal2 ;
        RECT 687.310 22.805 687.625 33.490 ;
        RECT 690.635 25.675 691.015 26.055 ;
        RECT 692.700 25.650 693.010 29.770 ;
        RECT 705.770 29.345 706.065 34.715 ;
      LAYER Metal3 ;
        RECT 705.770 34.260 721.790 34.670 ;
        RECT 690.635 25.665 693.115 26.065 ;
    END
  END b4_r7_b
  PIN b5_r0_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 864.060 171.120 865.260 171.500 ;
        RECT 864.060 168.820 867.320 169.200 ;
        RECT 864.725 166.905 887.280 167.245 ;
        RECT 888.390 166.915 903.035 167.215 ;
        RECT 864.040 163.320 867.340 163.700 ;
        RECT 891.415 163.240 894.335 163.540 ;
        RECT 897.880 163.225 901.250 163.525 ;
        RECT 864.040 161.320 865.325 161.700 ;
      LAYER Metal2 ;
        RECT 864.885 160.590 865.200 171.640 ;
        RECT 886.860 166.835 887.280 167.295 ;
        RECT 888.360 166.830 888.780 167.290 ;
        RECT 891.450 163.190 891.750 167.250 ;
        RECT 897.940 163.175 898.220 167.265 ;
        RECT 902.705 166.785 903.010 172.260 ;
      LAYER Metal3 ;
        RECT 902.660 171.750 918.140 172.205 ;
        RECT 886.830 166.885 888.855 167.270 ;
    END
  END b5_r0_b_not
  PIN b5_r1_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 863.860 151.395 865.060 151.775 ;
        RECT 863.860 149.095 867.120 149.475 ;
        RECT 864.525 147.180 887.080 147.520 ;
        RECT 888.190 147.190 902.835 147.490 ;
        RECT 863.840 143.595 867.140 143.975 ;
        RECT 891.215 143.515 894.135 143.815 ;
        RECT 897.680 143.500 901.050 143.800 ;
        RECT 863.840 141.595 865.125 141.975 ;
      LAYER Metal2 ;
        RECT 864.685 140.865 865.000 151.915 ;
        RECT 886.660 147.110 887.080 147.570 ;
        RECT 888.160 147.105 888.580 147.565 ;
        RECT 891.250 143.465 891.550 147.525 ;
        RECT 897.740 143.450 898.020 147.540 ;
        RECT 902.505 147.060 902.810 152.535 ;
      LAYER Metal3 ;
        RECT 902.460 152.025 917.940 152.480 ;
        RECT 886.630 147.160 888.655 147.545 ;
    END
  END b5_r1_b_not
  PIN b5_r0_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 883.585 171.220 884.820 171.600 ;
        RECT 881.560 168.820 884.820 169.200 ;
        RECT 888.990 167.660 902.605 167.960 ;
        RECT 890.185 165.005 894.315 165.305 ;
        RECT 896.690 164.955 901.190 165.265 ;
        RECT 883.445 163.960 887.390 164.295 ;
        RECT 881.540 163.320 884.840 163.700 ;
        RECT 883.355 161.320 884.840 161.700 ;
      LAYER Metal2 ;
        RECT 883.670 161.075 883.985 171.760 ;
        RECT 886.995 163.945 887.375 164.325 ;
        RECT 889.060 163.920 889.370 168.040 ;
        RECT 902.130 167.615 902.425 172.985 ;
      LAYER Metal3 ;
        RECT 902.130 172.530 918.150 172.940 ;
        RECT 886.995 163.935 889.475 164.335 ;
    END
  END b5_r0_b
  PIN b5_r1_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 883.385 151.495 884.620 151.875 ;
        RECT 881.360 149.095 884.620 149.475 ;
        RECT 888.790 147.935 902.405 148.235 ;
        RECT 889.985 145.280 894.115 145.580 ;
        RECT 896.490 145.230 900.990 145.540 ;
        RECT 883.245 144.235 887.190 144.570 ;
        RECT 881.340 143.595 884.640 143.975 ;
        RECT 883.155 141.595 884.640 141.975 ;
      LAYER Metal2 ;
        RECT 883.470 141.350 883.785 152.035 ;
        RECT 886.795 144.220 887.175 144.600 ;
        RECT 888.860 144.195 889.170 148.315 ;
        RECT 901.930 147.890 902.225 153.260 ;
      LAYER Metal3 ;
        RECT 901.930 152.805 917.950 153.215 ;
        RECT 886.795 144.210 889.275 144.610 ;
    END
  END b5_r1_b
  PIN b5_r2_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 864.015 131.750 865.215 132.130 ;
        RECT 864.015 129.450 867.275 129.830 ;
        RECT 864.680 127.535 887.235 127.875 ;
        RECT 888.345 127.545 902.990 127.845 ;
        RECT 863.995 123.950 867.295 124.330 ;
        RECT 891.370 123.870 894.290 124.170 ;
        RECT 897.835 123.855 901.205 124.155 ;
        RECT 863.995 121.950 865.280 122.330 ;
      LAYER Metal2 ;
        RECT 864.840 121.220 865.155 132.270 ;
        RECT 886.815 127.465 887.235 127.925 ;
        RECT 888.315 127.460 888.735 127.920 ;
        RECT 891.405 123.820 891.705 127.880 ;
        RECT 897.895 123.805 898.175 127.895 ;
        RECT 902.660 127.415 902.965 132.890 ;
      LAYER Metal3 ;
        RECT 902.615 132.380 918.095 132.835 ;
        RECT 886.785 127.515 888.810 127.900 ;
    END
  END b5_r2_b_not
  PIN b5_r2_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 883.540 131.850 884.775 132.230 ;
        RECT 881.515 129.450 884.775 129.830 ;
        RECT 888.945 128.290 902.560 128.590 ;
        RECT 890.140 125.635 894.270 125.935 ;
        RECT 896.645 125.585 901.145 125.895 ;
        RECT 883.400 124.590 887.345 124.925 ;
        RECT 881.495 123.950 884.795 124.330 ;
        RECT 883.310 121.950 884.795 122.330 ;
      LAYER Metal2 ;
        RECT 883.625 121.705 883.940 132.390 ;
        RECT 886.950 124.575 887.330 124.955 ;
        RECT 889.015 124.550 889.325 128.670 ;
        RECT 902.085 128.245 902.380 133.615 ;
      LAYER Metal3 ;
        RECT 902.085 133.160 918.105 133.570 ;
        RECT 886.950 124.565 889.430 124.965 ;
    END
  END b5_r2_b
  PIN b5_r3_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 864.015 111.955 865.215 112.335 ;
        RECT 864.015 109.655 867.275 110.035 ;
        RECT 864.680 107.740 887.235 108.080 ;
        RECT 888.345 107.750 902.990 108.050 ;
        RECT 863.995 104.155 867.295 104.535 ;
        RECT 891.370 104.075 894.290 104.375 ;
        RECT 897.835 104.060 901.205 104.360 ;
        RECT 863.995 102.155 865.280 102.535 ;
      LAYER Metal2 ;
        RECT 864.840 101.425 865.155 112.475 ;
        RECT 886.815 107.670 887.235 108.130 ;
        RECT 888.315 107.665 888.735 108.125 ;
        RECT 891.405 104.025 891.705 108.085 ;
        RECT 897.895 104.010 898.175 108.100 ;
        RECT 902.660 107.620 902.965 113.095 ;
      LAYER Metal3 ;
        RECT 902.615 112.585 918.095 113.040 ;
        RECT 886.785 107.720 888.810 108.105 ;
    END
  END b5_r3_b_not
  PIN b5_r3_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 883.540 112.055 884.775 112.435 ;
        RECT 881.515 109.655 884.775 110.035 ;
        RECT 888.945 108.495 902.560 108.795 ;
        RECT 890.140 105.840 894.270 106.140 ;
        RECT 896.645 105.790 901.145 106.100 ;
        RECT 883.400 104.795 887.345 105.130 ;
        RECT 881.495 104.155 884.795 104.535 ;
        RECT 883.310 102.155 884.795 102.535 ;
      LAYER Metal2 ;
        RECT 883.625 101.910 883.940 112.595 ;
        RECT 886.950 104.780 887.330 105.160 ;
        RECT 889.015 104.755 889.325 108.875 ;
        RECT 902.085 108.450 902.380 113.820 ;
      LAYER Metal3 ;
        RECT 902.085 113.365 918.105 113.775 ;
        RECT 886.950 104.770 889.430 105.170 ;
    END
  END b5_r3_b
  PIN b5_r4_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 863.935 92.200 865.135 92.580 ;
        RECT 863.935 89.900 867.195 90.280 ;
        RECT 864.600 87.985 887.155 88.325 ;
        RECT 888.265 87.995 902.910 88.295 ;
        RECT 863.915 84.400 867.215 84.780 ;
        RECT 891.290 84.320 894.210 84.620 ;
        RECT 897.755 84.305 901.125 84.605 ;
        RECT 863.915 82.400 865.200 82.780 ;
      LAYER Metal2 ;
        RECT 864.760 81.670 865.075 92.720 ;
        RECT 886.735 87.915 887.155 88.375 ;
        RECT 888.235 87.910 888.655 88.370 ;
        RECT 891.325 84.270 891.625 88.330 ;
        RECT 897.815 84.255 898.095 88.345 ;
        RECT 902.580 87.865 902.885 93.340 ;
      LAYER Metal3 ;
        RECT 902.535 92.830 918.015 93.285 ;
        RECT 886.705 87.965 888.730 88.350 ;
    END
  END b5_r4_b_not
  PIN b5_r4_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 883.460 92.300 884.695 92.680 ;
        RECT 881.435 89.900 884.695 90.280 ;
        RECT 888.865 88.740 902.480 89.040 ;
        RECT 890.060 86.085 894.190 86.385 ;
        RECT 896.565 86.035 901.065 86.345 ;
        RECT 883.320 85.040 887.265 85.375 ;
        RECT 881.415 84.400 884.715 84.780 ;
        RECT 883.230 82.400 884.715 82.780 ;
      LAYER Metal2 ;
        RECT 883.545 82.155 883.860 92.840 ;
        RECT 886.870 85.025 887.250 85.405 ;
        RECT 888.935 85.000 889.245 89.120 ;
        RECT 902.005 88.695 902.300 94.065 ;
      LAYER Metal3 ;
        RECT 902.005 93.610 918.025 94.020 ;
        RECT 886.870 85.015 889.350 85.415 ;
    END
  END b5_r4_b
  PIN b5_r5_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 864.040 72.485 865.240 72.865 ;
        RECT 864.040 70.185 867.300 70.565 ;
        RECT 864.705 68.270 887.260 68.610 ;
        RECT 888.370 68.280 903.015 68.580 ;
        RECT 864.020 64.685 867.320 65.065 ;
        RECT 891.395 64.605 894.315 64.905 ;
        RECT 897.860 64.590 901.230 64.890 ;
        RECT 864.020 62.685 865.305 63.065 ;
      LAYER Metal2 ;
        RECT 864.865 61.955 865.180 73.005 ;
        RECT 886.840 68.200 887.260 68.660 ;
        RECT 888.340 68.195 888.760 68.655 ;
        RECT 891.430 64.555 891.730 68.615 ;
        RECT 897.920 64.540 898.200 68.630 ;
        RECT 902.685 68.150 902.990 73.625 ;
      LAYER Metal3 ;
        RECT 902.640 73.115 918.120 73.570 ;
        RECT 886.810 68.250 888.835 68.635 ;
    END
  END b5_r5_b_not
  PIN b5_r5_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 883.565 72.585 884.800 72.965 ;
        RECT 881.540 70.185 884.800 70.565 ;
        RECT 888.970 69.025 902.585 69.325 ;
        RECT 890.165 66.370 894.295 66.670 ;
        RECT 896.670 66.320 901.170 66.630 ;
        RECT 883.425 65.325 887.370 65.660 ;
        RECT 881.520 64.685 884.820 65.065 ;
        RECT 883.335 62.685 884.820 63.065 ;
      LAYER Metal2 ;
        RECT 883.650 62.440 883.965 73.125 ;
        RECT 886.975 65.310 887.355 65.690 ;
        RECT 889.040 65.285 889.350 69.405 ;
        RECT 902.110 68.980 902.405 74.350 ;
      LAYER Metal3 ;
        RECT 902.110 73.895 918.130 74.305 ;
        RECT 886.975 65.300 889.455 65.700 ;
    END
  END b5_r5_b
  PIN b5_r6_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 864.040 52.515 865.240 52.895 ;
        RECT 864.040 50.215 867.300 50.595 ;
        RECT 864.705 48.300 887.260 48.640 ;
        RECT 888.370 48.310 903.015 48.610 ;
        RECT 864.020 44.715 867.320 45.095 ;
        RECT 891.395 44.635 894.315 44.935 ;
        RECT 897.860 44.620 901.230 44.920 ;
        RECT 864.020 42.715 865.305 43.095 ;
      LAYER Metal2 ;
        RECT 864.865 41.985 865.180 53.035 ;
        RECT 886.840 48.230 887.260 48.690 ;
        RECT 888.340 48.225 888.760 48.685 ;
        RECT 891.430 44.585 891.730 48.645 ;
        RECT 897.920 44.570 898.200 48.660 ;
        RECT 902.685 48.180 902.990 53.655 ;
      LAYER Metal3 ;
        RECT 902.640 53.145 918.120 53.600 ;
        RECT 886.810 48.280 888.835 48.665 ;
    END
  END b5_r6_b_not
  PIN b5_r6_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 883.565 52.615 884.800 52.995 ;
        RECT 881.540 50.215 884.800 50.595 ;
        RECT 888.970 49.055 902.585 49.355 ;
        RECT 890.165 46.400 894.295 46.700 ;
        RECT 896.670 46.350 901.170 46.660 ;
        RECT 883.425 45.355 887.370 45.690 ;
        RECT 881.520 44.715 884.820 45.095 ;
        RECT 883.335 42.715 884.820 43.095 ;
      LAYER Metal2 ;
        RECT 883.650 42.470 883.965 53.155 ;
        RECT 886.975 45.340 887.355 45.720 ;
        RECT 889.040 45.315 889.350 49.435 ;
        RECT 902.110 49.010 902.405 54.380 ;
      LAYER Metal3 ;
        RECT 902.110 53.925 918.130 54.335 ;
        RECT 886.975 45.330 889.455 45.730 ;
    END
  END b5_r6_b
  PIN b5_r7_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 864.040 32.850 865.240 33.230 ;
        RECT 864.040 30.550 867.300 30.930 ;
        RECT 864.705 28.635 887.260 28.975 ;
        RECT 888.370 28.645 903.015 28.945 ;
        RECT 864.020 25.050 867.320 25.430 ;
        RECT 891.395 24.970 894.315 25.270 ;
        RECT 897.860 24.955 901.230 25.255 ;
        RECT 864.020 23.050 865.305 23.430 ;
      LAYER Metal2 ;
        RECT 864.865 22.320 865.180 33.370 ;
        RECT 886.840 28.565 887.260 29.025 ;
        RECT 888.340 28.560 888.760 29.020 ;
        RECT 891.430 24.920 891.730 28.980 ;
        RECT 897.920 24.905 898.200 28.995 ;
        RECT 902.685 28.515 902.990 33.990 ;
      LAYER Metal3 ;
        RECT 902.640 33.480 918.120 33.935 ;
        RECT 886.810 28.615 888.835 29.000 ;
    END
  END b5_r7_b_not
  PIN b5_r7_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 883.565 32.950 884.800 33.330 ;
        RECT 881.540 30.550 884.800 30.930 ;
        RECT 888.970 29.390 902.585 29.690 ;
        RECT 890.165 26.735 894.295 27.035 ;
        RECT 896.670 26.685 901.170 26.995 ;
        RECT 883.425 25.690 887.370 26.025 ;
        RECT 881.520 25.050 884.820 25.430 ;
        RECT 883.335 23.050 884.820 23.430 ;
      LAYER Metal2 ;
        RECT 883.650 22.805 883.965 33.490 ;
        RECT 886.975 25.675 887.355 26.055 ;
        RECT 889.040 25.650 889.350 29.770 ;
        RECT 902.110 29.345 902.405 34.715 ;
      LAYER Metal3 ;
        RECT 902.110 34.260 918.130 34.670 ;
        RECT 886.975 25.665 889.455 26.065 ;
    END
  END b5_r7_b
  PIN b6_r0_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1060.400 171.120 1061.600 171.500 ;
        RECT 1060.400 168.820 1063.660 169.200 ;
        RECT 1061.065 166.905 1083.620 167.245 ;
        RECT 1084.730 166.915 1099.375 167.215 ;
        RECT 1060.380 163.320 1063.680 163.700 ;
        RECT 1087.755 163.240 1090.675 163.540 ;
        RECT 1094.220 163.225 1097.590 163.525 ;
        RECT 1060.380 161.320 1061.665 161.700 ;
      LAYER Metal2 ;
        RECT 1061.225 160.590 1061.540 171.640 ;
        RECT 1083.200 166.835 1083.620 167.295 ;
        RECT 1084.700 166.830 1085.120 167.290 ;
        RECT 1087.790 163.190 1088.090 167.250 ;
        RECT 1094.280 163.175 1094.560 167.265 ;
        RECT 1099.045 166.785 1099.350 172.260 ;
      LAYER Metal3 ;
        RECT 1099.000 171.750 1114.480 172.205 ;
        RECT 1083.170 166.885 1085.195 167.270 ;
    END
  END b6_r0_b_not
  PIN b6_r1_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1060.200 151.395 1061.400 151.775 ;
        RECT 1060.200 149.095 1063.460 149.475 ;
        RECT 1060.865 147.180 1083.420 147.520 ;
        RECT 1084.530 147.190 1099.175 147.490 ;
        RECT 1060.180 143.595 1063.480 143.975 ;
        RECT 1087.555 143.515 1090.475 143.815 ;
        RECT 1094.020 143.500 1097.390 143.800 ;
        RECT 1060.180 141.595 1061.465 141.975 ;
      LAYER Metal2 ;
        RECT 1061.025 140.865 1061.340 151.915 ;
        RECT 1083.000 147.110 1083.420 147.570 ;
        RECT 1084.500 147.105 1084.920 147.565 ;
        RECT 1087.590 143.465 1087.890 147.525 ;
        RECT 1094.080 143.450 1094.360 147.540 ;
        RECT 1098.845 147.060 1099.150 152.535 ;
      LAYER Metal3 ;
        RECT 1098.800 152.025 1114.280 152.480 ;
        RECT 1082.970 147.160 1084.995 147.545 ;
    END
  END b6_r1_b_not
  PIN b6_r0_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1079.925 171.220 1081.160 171.600 ;
        RECT 1077.900 168.820 1081.160 169.200 ;
        RECT 1085.330 167.660 1098.945 167.960 ;
        RECT 1086.525 165.005 1090.655 165.305 ;
        RECT 1093.030 164.955 1097.530 165.265 ;
        RECT 1079.785 163.960 1083.730 164.295 ;
        RECT 1077.880 163.320 1081.180 163.700 ;
        RECT 1079.695 161.320 1081.180 161.700 ;
      LAYER Metal2 ;
        RECT 1080.010 161.075 1080.325 171.760 ;
        RECT 1083.335 163.945 1083.715 164.325 ;
        RECT 1085.400 163.920 1085.710 168.040 ;
        RECT 1098.470 167.615 1098.765 172.985 ;
      LAYER Metal3 ;
        RECT 1098.470 172.530 1114.490 172.940 ;
        RECT 1083.335 163.935 1085.815 164.335 ;
    END
  END b6_r0_b
  PIN b6_r1_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1079.725 151.495 1080.960 151.875 ;
        RECT 1077.700 149.095 1080.960 149.475 ;
        RECT 1085.130 147.935 1098.745 148.235 ;
        RECT 1086.325 145.280 1090.455 145.580 ;
        RECT 1092.830 145.230 1097.330 145.540 ;
        RECT 1079.585 144.235 1083.530 144.570 ;
        RECT 1077.680 143.595 1080.980 143.975 ;
        RECT 1079.495 141.595 1080.980 141.975 ;
      LAYER Metal2 ;
        RECT 1079.810 141.350 1080.125 152.035 ;
        RECT 1083.135 144.220 1083.515 144.600 ;
        RECT 1085.200 144.195 1085.510 148.315 ;
        RECT 1098.270 147.890 1098.565 153.260 ;
      LAYER Metal3 ;
        RECT 1098.270 152.805 1114.290 153.215 ;
        RECT 1083.135 144.210 1085.615 144.610 ;
    END
  END b6_r1_b
  PIN b6_r2_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1060.355 131.750 1061.555 132.130 ;
        RECT 1060.355 129.450 1063.615 129.830 ;
        RECT 1061.020 127.535 1083.575 127.875 ;
        RECT 1084.685 127.545 1099.330 127.845 ;
        RECT 1060.335 123.950 1063.635 124.330 ;
        RECT 1087.710 123.870 1090.630 124.170 ;
        RECT 1094.175 123.855 1097.545 124.155 ;
        RECT 1060.335 121.950 1061.620 122.330 ;
      LAYER Metal2 ;
        RECT 1061.180 121.220 1061.495 132.270 ;
        RECT 1083.155 127.465 1083.575 127.925 ;
        RECT 1084.655 127.460 1085.075 127.920 ;
        RECT 1087.745 123.820 1088.045 127.880 ;
        RECT 1094.235 123.805 1094.515 127.895 ;
        RECT 1099.000 127.415 1099.305 132.890 ;
      LAYER Metal3 ;
        RECT 1098.955 132.380 1114.435 132.835 ;
        RECT 1083.125 127.515 1085.150 127.900 ;
    END
  END b6_r2_b_not
  PIN b6_r2_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1079.880 131.850 1081.115 132.230 ;
        RECT 1077.855 129.450 1081.115 129.830 ;
        RECT 1085.285 128.290 1098.900 128.590 ;
        RECT 1086.480 125.635 1090.610 125.935 ;
        RECT 1092.985 125.585 1097.485 125.895 ;
        RECT 1079.740 124.590 1083.685 124.925 ;
        RECT 1077.835 123.950 1081.135 124.330 ;
        RECT 1079.650 121.950 1081.135 122.330 ;
      LAYER Metal2 ;
        RECT 1079.965 121.705 1080.280 132.390 ;
        RECT 1083.290 124.575 1083.670 124.955 ;
        RECT 1085.355 124.550 1085.665 128.670 ;
        RECT 1098.425 128.245 1098.720 133.615 ;
      LAYER Metal3 ;
        RECT 1098.425 133.160 1114.445 133.570 ;
        RECT 1083.290 124.565 1085.770 124.965 ;
    END
  END b6_r2_b
  PIN b6_r3_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1060.355 111.955 1061.555 112.335 ;
        RECT 1060.355 109.655 1063.615 110.035 ;
        RECT 1061.020 107.740 1083.575 108.080 ;
        RECT 1084.685 107.750 1099.330 108.050 ;
        RECT 1060.335 104.155 1063.635 104.535 ;
        RECT 1087.710 104.075 1090.630 104.375 ;
        RECT 1094.175 104.060 1097.545 104.360 ;
        RECT 1060.335 102.155 1061.620 102.535 ;
      LAYER Metal2 ;
        RECT 1061.180 101.425 1061.495 112.475 ;
        RECT 1083.155 107.670 1083.575 108.130 ;
        RECT 1084.655 107.665 1085.075 108.125 ;
        RECT 1087.745 104.025 1088.045 108.085 ;
        RECT 1094.235 104.010 1094.515 108.100 ;
        RECT 1099.000 107.620 1099.305 113.095 ;
      LAYER Metal3 ;
        RECT 1098.955 112.585 1114.435 113.040 ;
        RECT 1083.125 107.720 1085.150 108.105 ;
    END
  END b6_r3_b_not
  PIN b6_r3_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1079.880 112.055 1081.115 112.435 ;
        RECT 1077.855 109.655 1081.115 110.035 ;
        RECT 1085.285 108.495 1098.900 108.795 ;
        RECT 1086.480 105.840 1090.610 106.140 ;
        RECT 1092.985 105.790 1097.485 106.100 ;
        RECT 1079.740 104.795 1083.685 105.130 ;
        RECT 1077.835 104.155 1081.135 104.535 ;
        RECT 1079.650 102.155 1081.135 102.535 ;
      LAYER Metal2 ;
        RECT 1079.965 101.910 1080.280 112.595 ;
        RECT 1083.290 104.780 1083.670 105.160 ;
        RECT 1085.355 104.755 1085.665 108.875 ;
        RECT 1098.425 108.450 1098.720 113.820 ;
      LAYER Metal3 ;
        RECT 1098.425 113.365 1114.445 113.775 ;
        RECT 1083.290 104.770 1085.770 105.170 ;
    END
  END b6_r3_b
  PIN b6_r4_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1060.275 92.200 1061.475 92.580 ;
        RECT 1060.275 89.900 1063.535 90.280 ;
        RECT 1060.940 87.985 1083.495 88.325 ;
        RECT 1084.605 87.995 1099.250 88.295 ;
        RECT 1060.255 84.400 1063.555 84.780 ;
        RECT 1087.630 84.320 1090.550 84.620 ;
        RECT 1094.095 84.305 1097.465 84.605 ;
        RECT 1060.255 82.400 1061.540 82.780 ;
      LAYER Metal2 ;
        RECT 1061.100 81.670 1061.415 92.720 ;
        RECT 1083.075 87.915 1083.495 88.375 ;
        RECT 1084.575 87.910 1084.995 88.370 ;
        RECT 1087.665 84.270 1087.965 88.330 ;
        RECT 1094.155 84.255 1094.435 88.345 ;
        RECT 1098.920 87.865 1099.225 93.340 ;
      LAYER Metal3 ;
        RECT 1098.875 92.830 1114.355 93.285 ;
        RECT 1083.045 87.965 1085.070 88.350 ;
    END
  END b6_r4_b_not
  PIN b6_r4_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1079.800 92.300 1081.035 92.680 ;
        RECT 1077.775 89.900 1081.035 90.280 ;
        RECT 1085.205 88.740 1098.820 89.040 ;
        RECT 1086.400 86.085 1090.530 86.385 ;
        RECT 1092.905 86.035 1097.405 86.345 ;
        RECT 1079.660 85.040 1083.605 85.375 ;
        RECT 1077.755 84.400 1081.055 84.780 ;
        RECT 1079.570 82.400 1081.055 82.780 ;
      LAYER Metal2 ;
        RECT 1079.885 82.155 1080.200 92.840 ;
        RECT 1083.210 85.025 1083.590 85.405 ;
        RECT 1085.275 85.000 1085.585 89.120 ;
        RECT 1098.345 88.695 1098.640 94.065 ;
      LAYER Metal3 ;
        RECT 1098.345 93.610 1114.365 94.020 ;
        RECT 1083.210 85.015 1085.690 85.415 ;
    END
  END b6_r4_b
  PIN b6_r5_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1060.380 72.485 1061.580 72.865 ;
        RECT 1060.380 70.185 1063.640 70.565 ;
        RECT 1061.045 68.270 1083.600 68.610 ;
        RECT 1084.710 68.280 1099.355 68.580 ;
        RECT 1060.360 64.685 1063.660 65.065 ;
        RECT 1087.735 64.605 1090.655 64.905 ;
        RECT 1094.200 64.590 1097.570 64.890 ;
        RECT 1060.360 62.685 1061.645 63.065 ;
      LAYER Metal2 ;
        RECT 1061.205 61.955 1061.520 73.005 ;
        RECT 1083.180 68.200 1083.600 68.660 ;
        RECT 1084.680 68.195 1085.100 68.655 ;
        RECT 1087.770 64.555 1088.070 68.615 ;
        RECT 1094.260 64.540 1094.540 68.630 ;
        RECT 1099.025 68.150 1099.330 73.625 ;
      LAYER Metal3 ;
        RECT 1098.980 73.115 1114.460 73.570 ;
        RECT 1083.150 68.250 1085.175 68.635 ;
    END
  END b6_r5_b_not
  PIN b6_r5_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1079.905 72.585 1081.140 72.965 ;
        RECT 1077.880 70.185 1081.140 70.565 ;
        RECT 1085.310 69.025 1098.925 69.325 ;
        RECT 1086.505 66.370 1090.635 66.670 ;
        RECT 1093.010 66.320 1097.510 66.630 ;
        RECT 1079.765 65.325 1083.710 65.660 ;
        RECT 1077.860 64.685 1081.160 65.065 ;
        RECT 1079.675 62.685 1081.160 63.065 ;
      LAYER Metal2 ;
        RECT 1079.990 62.440 1080.305 73.125 ;
        RECT 1083.315 65.310 1083.695 65.690 ;
        RECT 1085.380 65.285 1085.690 69.405 ;
        RECT 1098.450 68.980 1098.745 74.350 ;
      LAYER Metal3 ;
        RECT 1098.450 73.895 1114.470 74.305 ;
        RECT 1083.315 65.300 1085.795 65.700 ;
    END
  END b6_r5_b
  PIN b6_r6_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1060.380 52.515 1061.580 52.895 ;
        RECT 1060.380 50.215 1063.640 50.595 ;
        RECT 1061.045 48.300 1083.600 48.640 ;
        RECT 1084.710 48.310 1099.355 48.610 ;
        RECT 1060.360 44.715 1063.660 45.095 ;
        RECT 1087.735 44.635 1090.655 44.935 ;
        RECT 1094.200 44.620 1097.570 44.920 ;
        RECT 1060.360 42.715 1061.645 43.095 ;
      LAYER Metal2 ;
        RECT 1061.205 41.985 1061.520 53.035 ;
        RECT 1083.180 48.230 1083.600 48.690 ;
        RECT 1084.680 48.225 1085.100 48.685 ;
        RECT 1087.770 44.585 1088.070 48.645 ;
        RECT 1094.260 44.570 1094.540 48.660 ;
        RECT 1099.025 48.180 1099.330 53.655 ;
      LAYER Metal3 ;
        RECT 1098.980 53.145 1114.460 53.600 ;
        RECT 1083.150 48.280 1085.175 48.665 ;
    END
  END b6_r6_b_not
  PIN b6_r6_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1079.905 52.615 1081.140 52.995 ;
        RECT 1077.880 50.215 1081.140 50.595 ;
        RECT 1085.310 49.055 1098.925 49.355 ;
        RECT 1086.505 46.400 1090.635 46.700 ;
        RECT 1093.010 46.350 1097.510 46.660 ;
        RECT 1079.765 45.355 1083.710 45.690 ;
        RECT 1077.860 44.715 1081.160 45.095 ;
        RECT 1079.675 42.715 1081.160 43.095 ;
      LAYER Metal2 ;
        RECT 1079.990 42.470 1080.305 53.155 ;
        RECT 1083.315 45.340 1083.695 45.720 ;
        RECT 1085.380 45.315 1085.690 49.435 ;
        RECT 1098.450 49.010 1098.745 54.380 ;
      LAYER Metal3 ;
        RECT 1098.450 53.925 1114.470 54.335 ;
        RECT 1083.315 45.330 1085.795 45.730 ;
    END
  END b6_r6_b
  PIN b6_r7_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1060.380 32.850 1061.580 33.230 ;
        RECT 1060.380 30.550 1063.640 30.930 ;
        RECT 1061.045 28.635 1083.600 28.975 ;
        RECT 1084.710 28.645 1099.355 28.945 ;
        RECT 1060.360 25.050 1063.660 25.430 ;
        RECT 1087.735 24.970 1090.655 25.270 ;
        RECT 1094.200 24.955 1097.570 25.255 ;
        RECT 1060.360 23.050 1061.645 23.430 ;
      LAYER Metal2 ;
        RECT 1061.205 22.320 1061.520 33.370 ;
        RECT 1083.180 28.565 1083.600 29.025 ;
        RECT 1084.680 28.560 1085.100 29.020 ;
        RECT 1087.770 24.920 1088.070 28.980 ;
        RECT 1094.260 24.905 1094.540 28.995 ;
        RECT 1099.025 28.515 1099.330 33.990 ;
      LAYER Metal3 ;
        RECT 1098.980 33.480 1114.460 33.935 ;
        RECT 1083.150 28.615 1085.175 29.000 ;
    END
  END b6_r7_b_not
  PIN b6_r7_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 1079.905 32.950 1081.140 33.330 ;
        RECT 1077.880 30.550 1081.140 30.930 ;
        RECT 1085.310 29.390 1098.925 29.690 ;
        RECT 1086.505 26.735 1090.635 27.035 ;
        RECT 1093.010 26.685 1097.510 26.995 ;
        RECT 1079.765 25.690 1083.710 26.025 ;
        RECT 1077.860 25.050 1081.160 25.430 ;
        RECT 1079.675 23.050 1081.160 23.430 ;
      LAYER Metal2 ;
        RECT 1079.990 22.805 1080.305 33.490 ;
        RECT 1083.315 25.675 1083.695 26.055 ;
        RECT 1085.380 25.650 1085.690 29.770 ;
        RECT 1098.450 29.345 1098.745 34.715 ;
      LAYER Metal3 ;
        RECT 1098.450 34.260 1114.470 34.670 ;
        RECT 1083.315 25.665 1085.795 26.065 ;
    END
  END b6_r7_b
  PIN b0_r6_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 78.560 72.500 79.760 72.880 ;
        RECT 78.560 70.200 81.820 70.580 ;
        RECT 79.225 68.285 101.780 68.625 ;
        RECT 102.890 68.295 117.535 68.595 ;
        RECT 78.540 64.700 81.840 65.080 ;
        RECT 105.915 64.620 108.835 64.920 ;
        RECT 112.380 64.605 115.750 64.905 ;
        RECT 78.540 62.700 79.825 63.080 ;
      LAYER Metal2 ;
        RECT 79.385 61.970 79.700 73.020 ;
        RECT 101.360 68.215 101.780 68.675 ;
        RECT 102.860 68.210 103.280 68.670 ;
        RECT 105.950 64.570 106.250 68.630 ;
        RECT 112.440 64.555 112.720 68.645 ;
        RECT 117.205 68.165 117.510 73.640 ;
      LAYER Metal3 ;
        RECT 117.160 73.130 132.640 73.585 ;
        RECT 101.330 68.265 103.355 68.650 ;
    END
  END b0_r6_b_not
  PIN b3_r6_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 471.325 52.480 472.525 52.860 ;
        RECT 471.325 50.180 474.585 50.560 ;
        RECT 471.990 48.265 494.545 48.605 ;
        RECT 495.655 48.275 510.300 48.575 ;
        RECT 471.305 44.680 474.605 45.060 ;
        RECT 498.680 44.600 501.600 44.900 ;
        RECT 505.145 44.585 508.515 44.885 ;
        RECT 471.305 42.680 472.590 43.060 ;
      LAYER Metal2 ;
        RECT 472.150 41.950 472.465 53.000 ;
        RECT 494.125 48.195 494.545 48.655 ;
        RECT 495.625 48.190 496.045 48.650 ;
        RECT 498.715 44.550 499.015 48.610 ;
        RECT 505.205 44.535 505.485 48.625 ;
        RECT 509.970 48.145 510.275 53.620 ;
      LAYER Metal3 ;
        RECT 509.925 53.110 525.405 53.565 ;
        RECT 494.095 48.245 496.120 48.630 ;
    END
  END b3_r6_b_not
  PIN b3_r6_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 490.850 52.580 492.085 52.960 ;
        RECT 488.825 50.180 492.085 50.560 ;
        RECT 496.255 49.020 509.870 49.320 ;
        RECT 497.450 46.365 501.580 46.665 ;
        RECT 503.955 46.315 508.455 46.625 ;
        RECT 490.710 45.320 494.655 45.655 ;
        RECT 488.805 44.680 492.105 45.060 ;
        RECT 490.620 42.680 492.105 43.060 ;
      LAYER Metal2 ;
        RECT 490.935 42.435 491.250 53.120 ;
        RECT 494.260 45.305 494.640 45.685 ;
        RECT 496.325 45.280 496.635 49.400 ;
        RECT 509.395 48.975 509.690 54.345 ;
      LAYER Metal3 ;
        RECT 509.395 53.890 525.415 54.300 ;
        RECT 494.260 45.295 496.740 45.695 ;
    END
  END b3_r6_b
  PIN b3_r7_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 471.325 32.815 472.525 33.195 ;
        RECT 471.325 30.515 474.585 30.895 ;
        RECT 471.990 28.600 494.545 28.940 ;
        RECT 495.655 28.610 510.300 28.910 ;
        RECT 471.305 25.015 474.605 25.395 ;
        RECT 498.680 24.935 501.600 25.235 ;
        RECT 505.145 24.920 508.515 25.220 ;
        RECT 471.305 23.015 472.590 23.395 ;
      LAYER Metal2 ;
        RECT 472.150 22.285 472.465 33.335 ;
        RECT 494.125 28.530 494.545 28.990 ;
        RECT 495.625 28.525 496.045 28.985 ;
        RECT 498.715 24.885 499.015 28.945 ;
        RECT 505.205 24.870 505.485 28.960 ;
        RECT 509.970 28.480 510.275 33.955 ;
      LAYER Metal3 ;
        RECT 509.925 33.445 525.405 33.900 ;
        RECT 494.095 28.580 496.120 28.965 ;
    END
  END b3_r7_b_not
  PIN b3_r7_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 490.850 32.915 492.085 33.295 ;
        RECT 488.825 30.515 492.085 30.895 ;
        RECT 496.255 29.355 509.870 29.655 ;
        RECT 497.450 26.700 501.580 27.000 ;
        RECT 503.955 26.650 508.455 26.960 ;
        RECT 490.710 25.655 494.655 25.990 ;
        RECT 488.805 25.015 492.105 25.395 ;
        RECT 490.620 23.015 492.105 23.395 ;
      LAYER Metal2 ;
        RECT 490.935 22.770 491.250 33.455 ;
        RECT 494.260 25.640 494.640 26.020 ;
        RECT 496.325 25.615 496.635 29.735 ;
        RECT 509.395 29.310 509.690 34.680 ;
      LAYER Metal3 ;
        RECT 509.395 34.225 525.415 34.635 ;
        RECT 494.260 25.630 496.740 26.030 ;
    END
  END b3_r7_b
  PIN x0_a7_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 61.360 32.975 62.640 33.355 ;
        RECT 47.860 30.575 49.045 30.955 ;
        RECT 61.360 30.575 62.375 30.955 ;
        RECT 5.200 29.415 18.765 29.730 ;
        RECT 20.655 29.415 34.480 29.715 ;
        RECT 36.155 27.895 62.385 28.285 ;
        RECT 6.430 26.760 10.560 27.060 ;
        RECT 12.935 26.710 17.435 27.020 ;
        RECT 21.890 26.760 26.020 27.060 ;
        RECT 28.395 26.710 32.895 27.020 ;
        RECT 47.840 25.075 49.200 25.455 ;
        RECT 61.340 25.075 62.520 25.455 ;
        RECT 61.340 23.075 62.415 23.455 ;
      LAYER Metal2 ;
        RECT 5.205 29.370 5.585 29.750 ;
        RECT 18.370 29.370 18.750 29.750 ;
        RECT 20.640 29.370 21.020 29.775 ;
        RECT 34.105 29.370 34.465 31.200 ;
        RECT 36.285 27.850 36.700 31.200 ;
        RECT 48.480 30.940 48.790 30.970 ;
        RECT 48.480 24.840 48.795 30.940 ;
        RECT 61.980 22.845 62.310 33.540 ;
      LAYER Metal3 ;
        RECT 34.050 30.815 36.755 31.155 ;
        RECT -0.360 29.645 5.620 29.715 ;
        RECT -4.085 29.410 5.620 29.645 ;
        RECT -4.085 29.350 0.145 29.410 ;
        RECT 18.315 29.400 21.060 29.730 ;
    END
  END x0_a7_f
  PIN x0_a7_f_not
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 37.665 32.875 39.120 33.255 ;
        RECT 37.825 30.575 39.120 30.955 ;
        RECT 51.310 30.575 52.620 30.955 ;
        RECT 36.155 29.250 52.165 29.625 ;
        RECT 5.195 28.670 18.755 28.970 ;
        RECT 20.660 28.670 39.080 28.970 ;
        RECT 7.660 24.995 10.580 25.295 ;
        RECT 14.125 24.980 17.495 25.280 ;
        RECT 23.120 24.995 26.040 25.295 ;
        RECT 29.585 24.980 32.955 25.280 ;
        RECT 37.835 25.075 39.140 25.455 ;
        RECT 51.175 25.075 52.640 25.455 ;
        RECT 37.650 23.075 39.140 23.455 ;
      LAYER Metal2 ;
        RECT 5.195 28.620 5.575 29.000 ;
        RECT 7.695 24.945 7.995 29.005 ;
        RECT 14.185 24.930 14.465 29.020 ;
        RECT 18.375 28.620 18.755 29.000 ;
        RECT 20.645 28.620 21.025 29.025 ;
        RECT 23.155 24.945 23.455 29.005 ;
        RECT 29.645 24.930 29.925 29.020 ;
        RECT 37.955 23.020 38.310 33.325 ;
        RECT 38.620 28.625 38.965 29.680 ;
        RECT 51.465 24.795 51.795 30.990 ;
      LAYER Metal3 ;
        RECT -2.190 28.675 5.600 28.970 ;
        RECT -2.190 28.625 0.125 28.675 ;
        RECT 18.320 28.650 21.060 28.980 ;
    END
  END x0_a7_f_not
  PIN x0_c0_f
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 27.935 168.955 28.315 169.335 ;
        RECT 26.335 168.440 27.535 168.730 ;
        RECT 20.270 166.270 27.530 166.570 ;
        RECT 27.125 162.665 28.315 162.950 ;
        RECT 26.345 162.000 26.725 162.380 ;
      LAYER Metal2 ;
        RECT 20.290 164.500 20.610 166.630 ;
        RECT 26.385 161.990 26.685 168.800 ;
        RECT 27.175 162.585 27.485 168.775 ;
        RECT 27.970 162.515 28.270 169.345 ;
      LAYER Metal3 ;
        RECT -0.210 164.570 20.675 164.865 ;
    END
  END x0_c0_f
  PIN x0_c0_f_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT 21.475 169.115 24.880 169.555 ;
        RECT 33.255 168.505 33.635 168.885 ;
        RECT 20.825 165.735 24.910 166.005 ;
        RECT 24.485 164.475 30.875 164.765 ;
        RECT 21.465 162.560 21.845 162.940 ;
        RECT 30.465 161.835 33.645 162.155 ;
      LAYER Metal2 ;
        RECT 20.900 163.660 21.180 166.065 ;
        RECT 21.510 162.505 21.810 169.545 ;
        RECT 24.535 164.375 24.860 169.535 ;
        RECT 30.545 161.775 30.825 164.810 ;
        RECT 33.295 161.730 33.595 168.885 ;
      LAYER Metal3 ;
        RECT -0.210 163.705 21.260 164.000 ;
    END
  END x0_c0_f_not
  PIN x0_a7_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 98.085 32.965 99.320 33.345 ;
        RECT 96.060 30.565 99.320 30.945 ;
        RECT 103.490 29.405 117.105 29.705 ;
        RECT 104.685 26.750 108.815 27.050 ;
        RECT 111.190 26.700 115.690 27.010 ;
        RECT 97.945 25.705 101.890 26.040 ;
        RECT 96.040 25.065 99.340 25.445 ;
        RECT 97.855 23.065 99.340 23.445 ;
      LAYER Metal2 ;
        RECT 98.170 22.820 98.485 33.505 ;
        RECT 101.495 25.690 101.875 26.070 ;
        RECT 103.560 25.665 103.870 29.785 ;
        RECT 116.630 29.360 116.925 34.730 ;
      LAYER Metal3 ;
        RECT 116.630 34.275 132.650 34.685 ;
        RECT 101.495 25.680 103.975 26.080 ;
    END
  END x0_a7_b
  PIN x0_a7_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 78.560 32.865 79.760 33.245 ;
        RECT 78.560 30.565 81.820 30.945 ;
        RECT 79.225 28.650 101.780 28.990 ;
        RECT 102.890 28.660 117.535 28.960 ;
        RECT 78.540 25.065 81.840 25.445 ;
        RECT 105.915 24.985 108.835 25.285 ;
        RECT 112.380 24.970 115.750 25.270 ;
        RECT 78.540 23.065 79.825 23.445 ;
      LAYER Metal2 ;
        RECT 79.385 22.335 79.700 33.385 ;
        RECT 101.360 28.580 101.780 29.040 ;
        RECT 102.860 28.575 103.280 29.035 ;
        RECT 105.950 24.935 106.250 28.995 ;
        RECT 112.440 24.920 112.720 29.010 ;
        RECT 117.205 28.530 117.510 34.005 ;
      LAYER Metal3 ;
        RECT 117.160 33.495 132.640 33.950 ;
        RECT 101.330 28.630 103.355 29.015 ;
    END
  END x0_a7_b_not
  PIN b0_r7_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 98.085 52.630 99.320 53.010 ;
        RECT 96.060 50.230 99.320 50.610 ;
        RECT 103.490 49.070 117.105 49.370 ;
        RECT 104.685 46.415 108.815 46.715 ;
        RECT 111.190 46.365 115.690 46.675 ;
        RECT 97.945 45.370 101.890 45.705 ;
        RECT 96.040 44.730 99.340 45.110 ;
        RECT 97.855 42.730 99.340 43.110 ;
      LAYER Metal2 ;
        RECT 98.170 42.485 98.485 53.170 ;
        RECT 101.495 45.355 101.875 45.735 ;
        RECT 103.560 45.330 103.870 49.450 ;
        RECT 116.630 49.025 116.925 54.395 ;
      LAYER Metal3 ;
        RECT 116.630 53.940 132.650 54.350 ;
        RECT 101.495 45.345 103.975 45.745 ;
    END
  END b0_r7_b
  PIN b0_r7_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 78.560 52.530 79.760 52.910 ;
        RECT 78.560 50.230 81.820 50.610 ;
        RECT 79.225 48.315 101.780 48.655 ;
        RECT 102.890 48.325 117.535 48.625 ;
        RECT 78.540 44.730 81.840 45.110 ;
        RECT 105.915 44.650 108.835 44.950 ;
        RECT 112.380 44.635 115.750 44.935 ;
        RECT 78.540 42.730 79.825 43.110 ;
      LAYER Metal2 ;
        RECT 79.385 42.000 79.700 53.050 ;
        RECT 101.360 48.245 101.780 48.705 ;
        RECT 102.860 48.240 103.280 48.700 ;
        RECT 105.950 44.600 106.250 48.660 ;
        RECT 112.440 44.585 112.720 48.675 ;
        RECT 117.205 48.195 117.510 53.670 ;
      LAYER Metal3 ;
        RECT 117.160 53.160 132.640 53.615 ;
        RECT 101.330 48.295 103.355 48.680 ;
    END
  END b0_r7_b_not
  PIN b0_r6_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 98.085 72.600 99.320 72.980 ;
        RECT 96.060 70.200 99.320 70.580 ;
        RECT 103.490 69.040 117.105 69.340 ;
        RECT 104.685 66.385 108.815 66.685 ;
        RECT 111.190 66.335 115.690 66.645 ;
        RECT 97.945 65.340 101.890 65.675 ;
        RECT 96.040 64.700 99.340 65.080 ;
        RECT 97.855 62.700 99.340 63.080 ;
      LAYER Metal2 ;
        RECT 98.170 62.455 98.485 73.140 ;
        RECT 101.495 65.325 101.875 65.705 ;
        RECT 103.560 65.300 103.870 69.420 ;
        RECT 116.630 68.995 116.925 74.365 ;
      LAYER Metal3 ;
        RECT 116.630 73.910 132.650 74.320 ;
        RECT 101.495 65.315 103.975 65.715 ;
    END
  END b0_r6_b
  PIN b0_r5_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 97.980 92.315 99.215 92.695 ;
        RECT 95.955 89.915 99.215 90.295 ;
        RECT 103.385 88.755 117.000 89.055 ;
        RECT 104.580 86.100 108.710 86.400 ;
        RECT 111.085 86.050 115.585 86.360 ;
        RECT 97.840 85.055 101.785 85.390 ;
        RECT 95.935 84.415 99.235 84.795 ;
        RECT 97.750 82.415 99.235 82.795 ;
      LAYER Metal2 ;
        RECT 98.065 82.170 98.380 92.855 ;
        RECT 101.390 85.040 101.770 85.420 ;
        RECT 103.455 85.015 103.765 89.135 ;
        RECT 116.525 88.710 116.820 94.080 ;
      LAYER Metal3 ;
        RECT 116.525 93.625 132.545 94.035 ;
        RECT 101.390 85.030 103.870 85.430 ;
    END
  END b0_r5_b
  PIN b0_r5_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 78.455 92.215 79.655 92.595 ;
        RECT 78.455 89.915 81.715 90.295 ;
        RECT 79.120 88.000 101.675 88.340 ;
        RECT 102.785 88.010 117.430 88.310 ;
        RECT 78.435 84.415 81.735 84.795 ;
        RECT 105.810 84.335 108.730 84.635 ;
        RECT 112.275 84.320 115.645 84.620 ;
        RECT 78.435 82.415 79.720 82.795 ;
      LAYER Metal2 ;
        RECT 79.280 81.685 79.595 92.735 ;
        RECT 101.255 87.930 101.675 88.390 ;
        RECT 102.755 87.925 103.175 88.385 ;
        RECT 105.845 84.285 106.145 88.345 ;
        RECT 112.335 84.270 112.615 88.360 ;
        RECT 117.100 87.880 117.405 93.355 ;
      LAYER Metal3 ;
        RECT 117.055 92.845 132.535 93.300 ;
        RECT 101.225 87.980 103.250 88.365 ;
    END
  END b0_r5_b_not
  PIN b0_r4_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 98.060 112.070 99.295 112.450 ;
        RECT 96.035 109.670 99.295 110.050 ;
        RECT 103.465 108.510 117.080 108.810 ;
        RECT 104.660 105.855 108.790 106.155 ;
        RECT 111.165 105.805 115.665 106.115 ;
        RECT 97.920 104.810 101.865 105.145 ;
        RECT 96.015 104.170 99.315 104.550 ;
        RECT 97.830 102.170 99.315 102.550 ;
      LAYER Metal2 ;
        RECT 98.145 101.925 98.460 112.610 ;
        RECT 101.470 104.795 101.850 105.175 ;
        RECT 103.535 104.770 103.845 108.890 ;
        RECT 116.605 108.465 116.900 113.835 ;
      LAYER Metal3 ;
        RECT 116.605 113.380 132.625 113.790 ;
        RECT 101.470 104.785 103.950 105.185 ;
    END
  END b0_r4_b
  PIN b0_r4_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 78.535 111.970 79.735 112.350 ;
        RECT 78.535 109.670 81.795 110.050 ;
        RECT 79.200 107.755 101.755 108.095 ;
        RECT 102.865 107.765 117.510 108.065 ;
        RECT 78.515 104.170 81.815 104.550 ;
        RECT 105.890 104.090 108.810 104.390 ;
        RECT 112.355 104.075 115.725 104.375 ;
        RECT 78.515 102.170 79.800 102.550 ;
      LAYER Metal2 ;
        RECT 79.360 101.440 79.675 112.490 ;
        RECT 101.335 107.685 101.755 108.145 ;
        RECT 102.835 107.680 103.255 108.140 ;
        RECT 105.925 104.040 106.225 108.100 ;
        RECT 112.415 104.025 112.695 108.115 ;
        RECT 117.180 107.635 117.485 113.110 ;
      LAYER Metal3 ;
        RECT 117.135 112.600 132.615 113.055 ;
        RECT 101.305 107.735 103.330 108.120 ;
    END
  END b0_r4_b_not
  PIN b0_r3_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 98.060 131.865 99.295 132.245 ;
        RECT 96.035 129.465 99.295 129.845 ;
        RECT 103.465 128.305 117.080 128.605 ;
        RECT 104.660 125.650 108.790 125.950 ;
        RECT 111.165 125.600 115.665 125.910 ;
        RECT 97.920 124.605 101.865 124.940 ;
        RECT 96.015 123.965 99.315 124.345 ;
        RECT 97.830 121.965 99.315 122.345 ;
      LAYER Metal2 ;
        RECT 98.145 121.720 98.460 132.405 ;
        RECT 101.470 124.590 101.850 124.970 ;
        RECT 103.535 124.565 103.845 128.685 ;
        RECT 116.605 128.260 116.900 133.630 ;
      LAYER Metal3 ;
        RECT 116.605 133.175 132.625 133.585 ;
        RECT 101.470 124.580 103.950 124.980 ;
    END
  END b0_r3_b
  PIN b0_r3_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 78.535 131.765 79.735 132.145 ;
        RECT 78.535 129.465 81.795 129.845 ;
        RECT 79.200 127.550 101.755 127.890 ;
        RECT 102.865 127.560 117.510 127.860 ;
        RECT 78.515 123.965 81.815 124.345 ;
        RECT 105.890 123.885 108.810 124.185 ;
        RECT 112.355 123.870 115.725 124.170 ;
        RECT 78.515 121.965 79.800 122.345 ;
      LAYER Metal2 ;
        RECT 79.360 121.235 79.675 132.285 ;
        RECT 101.335 127.480 101.755 127.940 ;
        RECT 102.835 127.475 103.255 127.935 ;
        RECT 105.925 123.835 106.225 127.895 ;
        RECT 112.415 123.820 112.695 127.910 ;
        RECT 117.180 127.430 117.485 132.905 ;
      LAYER Metal3 ;
        RECT 117.135 132.395 132.615 132.850 ;
        RECT 101.305 127.530 103.330 127.915 ;
    END
  END b0_r3_b_not
  PIN b0_r2_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 97.905 151.510 99.140 151.890 ;
        RECT 95.880 149.110 99.140 149.490 ;
        RECT 103.310 147.950 116.925 148.250 ;
        RECT 104.505 145.295 108.635 145.595 ;
        RECT 111.010 145.245 115.510 145.555 ;
        RECT 97.765 144.250 101.710 144.585 ;
        RECT 95.860 143.610 99.160 143.990 ;
        RECT 97.675 141.610 99.160 141.990 ;
      LAYER Metal2 ;
        RECT 97.990 141.365 98.305 152.050 ;
        RECT 101.315 144.235 101.695 144.615 ;
        RECT 103.380 144.210 103.690 148.330 ;
        RECT 116.450 147.905 116.745 153.275 ;
      LAYER Metal3 ;
        RECT 116.450 152.820 132.470 153.230 ;
        RECT 101.315 144.225 103.795 144.625 ;
    END
  END b0_r2_b
  PIN b0_r2_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 78.380 151.410 79.580 151.790 ;
        RECT 78.380 149.110 81.640 149.490 ;
        RECT 79.045 147.195 101.600 147.535 ;
        RECT 102.710 147.205 117.355 147.505 ;
        RECT 78.360 143.610 81.660 143.990 ;
        RECT 105.735 143.530 108.655 143.830 ;
        RECT 112.200 143.515 115.570 143.815 ;
        RECT 78.360 141.610 79.645 141.990 ;
      LAYER Metal2 ;
        RECT 79.205 140.880 79.520 151.930 ;
        RECT 101.180 147.125 101.600 147.585 ;
        RECT 102.680 147.120 103.100 147.580 ;
        RECT 105.770 143.480 106.070 147.540 ;
        RECT 112.260 143.465 112.540 147.555 ;
        RECT 117.025 147.075 117.330 152.550 ;
      LAYER Metal3 ;
        RECT 116.980 152.040 132.460 152.495 ;
        RECT 101.150 147.175 103.175 147.560 ;
    END
  END b0_r2_b_not
  PIN b0_r1_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 78.580 171.135 79.780 171.515 ;
        RECT 78.580 168.835 81.840 169.215 ;
        RECT 79.245 166.920 101.800 167.260 ;
        RECT 102.910 166.930 117.555 167.230 ;
        RECT 78.560 163.335 81.860 163.715 ;
        RECT 105.935 163.255 108.855 163.555 ;
        RECT 112.400 163.240 115.770 163.540 ;
        RECT 78.560 161.335 79.845 161.715 ;
      LAYER Metal2 ;
        RECT 79.405 160.605 79.720 171.655 ;
        RECT 101.380 166.850 101.800 167.310 ;
        RECT 102.880 166.845 103.300 167.305 ;
        RECT 105.970 163.205 106.270 167.265 ;
        RECT 112.460 163.190 112.740 167.280 ;
        RECT 117.225 166.800 117.530 172.275 ;
      LAYER Metal3 ;
        RECT 117.180 171.765 132.660 172.220 ;
        RECT 101.350 166.900 103.375 167.285 ;
    END
  END b0_r1_b_not
  PIN b0_r1_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 98.105 171.235 99.340 171.615 ;
        RECT 96.080 168.835 99.340 169.215 ;
        RECT 103.510 167.675 117.125 167.975 ;
        RECT 104.705 165.020 108.835 165.320 ;
        RECT 111.210 164.970 115.710 165.280 ;
        RECT 97.965 163.975 101.910 164.310 ;
        RECT 96.060 163.335 99.360 163.715 ;
        RECT 97.875 161.335 99.360 161.715 ;
      LAYER Metal2 ;
        RECT 98.190 161.090 98.505 171.775 ;
        RECT 101.515 163.960 101.895 164.340 ;
        RECT 103.580 163.935 103.890 168.055 ;
        RECT 116.650 167.630 116.945 173.000 ;
      LAYER Metal3 ;
        RECT 116.650 172.545 132.670 172.955 ;
        RECT 101.515 163.950 103.995 164.350 ;
    END
  END b0_r1_b
  PIN b2_r0_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 274.945 171.135 276.145 171.515 ;
        RECT 274.945 168.835 278.205 169.215 ;
        RECT 275.610 166.920 298.165 167.260 ;
        RECT 299.275 166.930 313.920 167.230 ;
        RECT 274.925 163.335 278.225 163.715 ;
        RECT 302.300 163.255 305.220 163.555 ;
        RECT 308.765 163.240 312.135 163.540 ;
        RECT 274.925 161.335 276.210 161.715 ;
      LAYER Metal2 ;
        RECT 275.770 160.605 276.085 171.655 ;
        RECT 297.745 166.850 298.165 167.310 ;
        RECT 299.245 166.845 299.665 167.305 ;
        RECT 302.335 163.205 302.635 167.265 ;
        RECT 308.825 163.190 309.105 167.280 ;
        RECT 313.590 166.800 313.895 172.275 ;
      LAYER Metal3 ;
        RECT 313.545 171.765 329.025 172.220 ;
        RECT 297.715 166.900 299.740 167.285 ;
    END
  END b2_r0_b_not
  PIN b2_r1_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 274.745 151.410 275.945 151.790 ;
        RECT 274.745 149.110 278.005 149.490 ;
        RECT 275.410 147.195 297.965 147.535 ;
        RECT 299.075 147.205 313.720 147.505 ;
        RECT 274.725 143.610 278.025 143.990 ;
        RECT 302.100 143.530 305.020 143.830 ;
        RECT 308.565 143.515 311.935 143.815 ;
        RECT 274.725 141.610 276.010 141.990 ;
      LAYER Metal2 ;
        RECT 275.570 140.880 275.885 151.930 ;
        RECT 297.545 147.125 297.965 147.585 ;
        RECT 299.045 147.120 299.465 147.580 ;
        RECT 302.135 143.480 302.435 147.540 ;
        RECT 308.625 143.465 308.905 147.555 ;
        RECT 313.390 147.075 313.695 152.550 ;
      LAYER Metal3 ;
        RECT 313.345 152.040 328.825 152.495 ;
        RECT 297.515 147.175 299.540 147.560 ;
    END
  END b2_r1_b_not
  PIN b2_r0_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 294.470 171.235 295.705 171.615 ;
        RECT 292.445 168.835 295.705 169.215 ;
        RECT 299.875 167.675 313.490 167.975 ;
        RECT 301.070 165.020 305.200 165.320 ;
        RECT 307.575 164.970 312.075 165.280 ;
        RECT 294.330 163.975 298.275 164.310 ;
        RECT 292.425 163.335 295.725 163.715 ;
        RECT 294.240 161.335 295.725 161.715 ;
      LAYER Metal2 ;
        RECT 294.555 161.090 294.870 171.775 ;
        RECT 297.880 163.960 298.260 164.340 ;
        RECT 299.945 163.935 300.255 168.055 ;
        RECT 313.015 167.630 313.310 173.000 ;
      LAYER Metal3 ;
        RECT 313.015 172.545 329.035 172.955 ;
        RECT 297.880 163.950 300.360 164.350 ;
    END
  END b2_r0_b
  PIN b2_r1_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 294.270 151.510 295.505 151.890 ;
        RECT 292.245 149.110 295.505 149.490 ;
        RECT 299.675 147.950 313.290 148.250 ;
        RECT 300.870 145.295 305.000 145.595 ;
        RECT 307.375 145.245 311.875 145.555 ;
        RECT 294.130 144.250 298.075 144.585 ;
        RECT 292.225 143.610 295.525 143.990 ;
        RECT 294.040 141.610 295.525 141.990 ;
      LAYER Metal2 ;
        RECT 294.355 141.365 294.670 152.050 ;
        RECT 297.680 144.235 298.060 144.615 ;
        RECT 299.745 144.210 300.055 148.330 ;
        RECT 312.815 147.905 313.110 153.275 ;
      LAYER Metal3 ;
        RECT 312.815 152.820 328.835 153.230 ;
        RECT 297.680 144.225 300.160 144.625 ;
    END
  END b2_r1_b
  PIN b2_r2_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 274.900 131.765 276.100 132.145 ;
        RECT 274.900 129.465 278.160 129.845 ;
        RECT 275.565 127.550 298.120 127.890 ;
        RECT 299.230 127.560 313.875 127.860 ;
        RECT 274.880 123.965 278.180 124.345 ;
        RECT 302.255 123.885 305.175 124.185 ;
        RECT 308.720 123.870 312.090 124.170 ;
        RECT 274.880 121.965 276.165 122.345 ;
      LAYER Metal2 ;
        RECT 275.725 121.235 276.040 132.285 ;
        RECT 297.700 127.480 298.120 127.940 ;
        RECT 299.200 127.475 299.620 127.935 ;
        RECT 302.290 123.835 302.590 127.895 ;
        RECT 308.780 123.820 309.060 127.910 ;
        RECT 313.545 127.430 313.850 132.905 ;
      LAYER Metal3 ;
        RECT 313.500 132.395 328.980 132.850 ;
        RECT 297.670 127.530 299.695 127.915 ;
    END
  END b2_r2_b_not
  PIN b2_r2_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 294.425 131.865 295.660 132.245 ;
        RECT 292.400 129.465 295.660 129.845 ;
        RECT 299.830 128.305 313.445 128.605 ;
        RECT 301.025 125.650 305.155 125.950 ;
        RECT 307.530 125.600 312.030 125.910 ;
        RECT 294.285 124.605 298.230 124.940 ;
        RECT 292.380 123.965 295.680 124.345 ;
        RECT 294.195 121.965 295.680 122.345 ;
      LAYER Metal2 ;
        RECT 294.510 121.720 294.825 132.405 ;
        RECT 297.835 124.590 298.215 124.970 ;
        RECT 299.900 124.565 300.210 128.685 ;
        RECT 312.970 128.260 313.265 133.630 ;
      LAYER Metal3 ;
        RECT 312.970 133.175 328.990 133.585 ;
        RECT 297.835 124.580 300.315 124.980 ;
    END
  END b2_r2_b
  PIN b2_r3_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 274.900 111.970 276.100 112.350 ;
        RECT 274.900 109.670 278.160 110.050 ;
        RECT 275.565 107.755 298.120 108.095 ;
        RECT 299.230 107.765 313.875 108.065 ;
        RECT 274.880 104.170 278.180 104.550 ;
        RECT 302.255 104.090 305.175 104.390 ;
        RECT 308.720 104.075 312.090 104.375 ;
        RECT 274.880 102.170 276.165 102.550 ;
      LAYER Metal2 ;
        RECT 275.725 101.440 276.040 112.490 ;
        RECT 297.700 107.685 298.120 108.145 ;
        RECT 299.200 107.680 299.620 108.140 ;
        RECT 302.290 104.040 302.590 108.100 ;
        RECT 308.780 104.025 309.060 108.115 ;
        RECT 313.545 107.635 313.850 113.110 ;
      LAYER Metal3 ;
        RECT 313.500 112.600 328.980 113.055 ;
        RECT 297.670 107.735 299.695 108.120 ;
    END
  END b2_r3_b_not
  PIN b2_r3_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 294.425 112.070 295.660 112.450 ;
        RECT 292.400 109.670 295.660 110.050 ;
        RECT 299.830 108.510 313.445 108.810 ;
        RECT 301.025 105.855 305.155 106.155 ;
        RECT 307.530 105.805 312.030 106.115 ;
        RECT 294.285 104.810 298.230 105.145 ;
        RECT 292.380 104.170 295.680 104.550 ;
        RECT 294.195 102.170 295.680 102.550 ;
      LAYER Metal2 ;
        RECT 294.510 101.925 294.825 112.610 ;
        RECT 297.835 104.795 298.215 105.175 ;
        RECT 299.900 104.770 300.210 108.890 ;
        RECT 312.970 108.465 313.265 113.835 ;
      LAYER Metal3 ;
        RECT 312.970 113.380 328.990 113.790 ;
        RECT 297.835 104.785 300.315 105.185 ;
    END
  END b2_r3_b
  PIN b2_r4_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 274.820 92.215 276.020 92.595 ;
        RECT 274.820 89.915 278.080 90.295 ;
        RECT 275.485 88.000 298.040 88.340 ;
        RECT 299.150 88.010 313.795 88.310 ;
        RECT 274.800 84.415 278.100 84.795 ;
        RECT 302.175 84.335 305.095 84.635 ;
        RECT 308.640 84.320 312.010 84.620 ;
        RECT 274.800 82.415 276.085 82.795 ;
      LAYER Metal2 ;
        RECT 275.645 81.685 275.960 92.735 ;
        RECT 297.620 87.930 298.040 88.390 ;
        RECT 299.120 87.925 299.540 88.385 ;
        RECT 302.210 84.285 302.510 88.345 ;
        RECT 308.700 84.270 308.980 88.360 ;
        RECT 313.465 87.880 313.770 93.355 ;
      LAYER Metal3 ;
        RECT 313.420 92.845 328.900 93.300 ;
        RECT 297.590 87.980 299.615 88.365 ;
    END
  END b2_r4_b_not
  PIN b2_r4_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 294.345 92.315 295.580 92.695 ;
        RECT 292.320 89.915 295.580 90.295 ;
        RECT 299.750 88.755 313.365 89.055 ;
        RECT 300.945 86.100 305.075 86.400 ;
        RECT 307.450 86.050 311.950 86.360 ;
        RECT 294.205 85.055 298.150 85.390 ;
        RECT 292.300 84.415 295.600 84.795 ;
        RECT 294.115 82.415 295.600 82.795 ;
      LAYER Metal2 ;
        RECT 294.430 82.170 294.745 92.855 ;
        RECT 297.755 85.040 298.135 85.420 ;
        RECT 299.820 85.015 300.130 89.135 ;
        RECT 312.890 88.710 313.185 94.080 ;
      LAYER Metal3 ;
        RECT 312.890 93.625 328.910 94.035 ;
        RECT 297.755 85.030 300.235 85.430 ;
    END
  END b2_r4_b
  PIN b2_r5_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 274.925 72.500 276.125 72.880 ;
        RECT 274.925 70.200 278.185 70.580 ;
        RECT 275.590 68.285 298.145 68.625 ;
        RECT 299.255 68.295 313.900 68.595 ;
        RECT 274.905 64.700 278.205 65.080 ;
        RECT 302.280 64.620 305.200 64.920 ;
        RECT 308.745 64.605 312.115 64.905 ;
        RECT 274.905 62.700 276.190 63.080 ;
      LAYER Metal2 ;
        RECT 275.750 61.970 276.065 73.020 ;
        RECT 297.725 68.215 298.145 68.675 ;
        RECT 299.225 68.210 299.645 68.670 ;
        RECT 302.315 64.570 302.615 68.630 ;
        RECT 308.805 64.555 309.085 68.645 ;
        RECT 313.570 68.165 313.875 73.640 ;
      LAYER Metal3 ;
        RECT 313.525 73.130 329.005 73.585 ;
        RECT 297.695 68.265 299.720 68.650 ;
    END
  END b2_r5_b_not
  PIN b2_r5_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 294.450 72.600 295.685 72.980 ;
        RECT 292.425 70.200 295.685 70.580 ;
        RECT 299.855 69.040 313.470 69.340 ;
        RECT 301.050 66.385 305.180 66.685 ;
        RECT 307.555 66.335 312.055 66.645 ;
        RECT 294.310 65.340 298.255 65.675 ;
        RECT 292.405 64.700 295.705 65.080 ;
        RECT 294.220 62.700 295.705 63.080 ;
      LAYER Metal2 ;
        RECT 294.535 62.455 294.850 73.140 ;
        RECT 297.860 65.325 298.240 65.705 ;
        RECT 299.925 65.300 300.235 69.420 ;
        RECT 312.995 68.995 313.290 74.365 ;
      LAYER Metal3 ;
        RECT 312.995 73.910 329.015 74.320 ;
        RECT 297.860 65.315 300.340 65.715 ;
    END
  END b2_r5_b
  PIN b2_r6_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 274.925 52.530 276.125 52.910 ;
        RECT 274.925 50.230 278.185 50.610 ;
        RECT 275.590 48.315 298.145 48.655 ;
        RECT 299.255 48.325 313.900 48.625 ;
        RECT 274.905 44.730 278.205 45.110 ;
        RECT 302.280 44.650 305.200 44.950 ;
        RECT 308.745 44.635 312.115 44.935 ;
        RECT 274.905 42.730 276.190 43.110 ;
      LAYER Metal2 ;
        RECT 275.750 42.000 276.065 53.050 ;
        RECT 297.725 48.245 298.145 48.705 ;
        RECT 299.225 48.240 299.645 48.700 ;
        RECT 302.315 44.600 302.615 48.660 ;
        RECT 308.805 44.585 309.085 48.675 ;
        RECT 313.570 48.195 313.875 53.670 ;
      LAYER Metal3 ;
        RECT 313.525 53.160 329.005 53.615 ;
        RECT 297.695 48.295 299.720 48.680 ;
    END
  END b2_r6_b_not
  PIN b2_r6_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 294.450 52.630 295.685 53.010 ;
        RECT 292.425 50.230 295.685 50.610 ;
        RECT 299.855 49.070 313.470 49.370 ;
        RECT 301.050 46.415 305.180 46.715 ;
        RECT 307.555 46.365 312.055 46.675 ;
        RECT 294.310 45.370 298.255 45.705 ;
        RECT 292.405 44.730 295.705 45.110 ;
        RECT 294.220 42.730 295.705 43.110 ;
      LAYER Metal2 ;
        RECT 294.535 42.485 294.850 53.170 ;
        RECT 297.860 45.355 298.240 45.735 ;
        RECT 299.925 45.330 300.235 49.450 ;
        RECT 312.995 49.025 313.290 54.395 ;
      LAYER Metal3 ;
        RECT 312.995 53.940 329.015 54.350 ;
        RECT 297.860 45.345 300.340 45.745 ;
    END
  END b2_r6_b
  PIN b2_r7_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 274.925 32.865 276.125 33.245 ;
        RECT 274.925 30.565 278.185 30.945 ;
        RECT 275.590 28.650 298.145 28.990 ;
        RECT 299.255 28.660 313.900 28.960 ;
        RECT 274.905 25.065 278.205 25.445 ;
        RECT 302.280 24.985 305.200 25.285 ;
        RECT 308.745 24.970 312.115 25.270 ;
        RECT 274.905 23.065 276.190 23.445 ;
      LAYER Metal2 ;
        RECT 275.750 22.335 276.065 33.385 ;
        RECT 297.725 28.580 298.145 29.040 ;
        RECT 299.225 28.575 299.645 29.035 ;
        RECT 302.315 24.935 302.615 28.995 ;
        RECT 308.805 24.920 309.085 29.010 ;
        RECT 313.570 28.530 313.875 34.005 ;
      LAYER Metal3 ;
        RECT 313.525 33.495 329.005 33.950 ;
        RECT 297.695 28.630 299.720 29.015 ;
    END
  END b2_r7_b_not
  PIN b2_r7_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 294.450 32.965 295.685 33.345 ;
        RECT 292.425 30.565 295.685 30.945 ;
        RECT 299.855 29.405 313.470 29.705 ;
        RECT 301.050 26.750 305.180 27.050 ;
        RECT 307.555 26.700 312.055 27.010 ;
        RECT 294.310 25.705 298.255 26.040 ;
        RECT 292.405 25.065 295.705 25.445 ;
        RECT 294.220 23.065 295.705 23.445 ;
      LAYER Metal2 ;
        RECT 294.535 22.820 294.850 33.505 ;
        RECT 297.860 25.690 298.240 26.070 ;
        RECT 299.925 25.665 300.235 29.785 ;
        RECT 312.995 29.360 313.290 34.730 ;
      LAYER Metal3 ;
        RECT 312.995 34.275 329.015 34.685 ;
        RECT 297.860 25.680 300.340 26.080 ;
    END
  END b2_r7_b
  PIN b3_r0_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 471.345 171.085 472.545 171.465 ;
        RECT 471.345 168.785 474.605 169.165 ;
        RECT 472.010 166.870 494.565 167.210 ;
        RECT 495.675 166.880 510.320 167.180 ;
        RECT 471.325 163.285 474.625 163.665 ;
        RECT 498.700 163.205 501.620 163.505 ;
        RECT 505.165 163.190 508.535 163.490 ;
        RECT 471.325 161.285 472.610 161.665 ;
      LAYER Metal2 ;
        RECT 472.170 160.555 472.485 171.605 ;
        RECT 494.145 166.800 494.565 167.260 ;
        RECT 495.645 166.795 496.065 167.255 ;
        RECT 498.735 163.155 499.035 167.215 ;
        RECT 505.225 163.140 505.505 167.230 ;
        RECT 509.990 166.750 510.295 172.225 ;
      LAYER Metal3 ;
        RECT 509.945 171.715 525.425 172.170 ;
        RECT 494.115 166.850 496.140 167.235 ;
    END
  END b3_r0_b_not
  PIN b3_r1_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 471.145 151.360 472.345 151.740 ;
        RECT 471.145 149.060 474.405 149.440 ;
        RECT 471.810 147.145 494.365 147.485 ;
        RECT 495.475 147.155 510.120 147.455 ;
        RECT 471.125 143.560 474.425 143.940 ;
        RECT 498.500 143.480 501.420 143.780 ;
        RECT 504.965 143.465 508.335 143.765 ;
        RECT 471.125 141.560 472.410 141.940 ;
      LAYER Metal2 ;
        RECT 471.970 140.830 472.285 151.880 ;
        RECT 493.945 147.075 494.365 147.535 ;
        RECT 495.445 147.070 495.865 147.530 ;
        RECT 498.535 143.430 498.835 147.490 ;
        RECT 505.025 143.415 505.305 147.505 ;
        RECT 509.790 147.025 510.095 152.500 ;
      LAYER Metal3 ;
        RECT 509.745 151.990 525.225 152.445 ;
        RECT 493.915 147.125 495.940 147.510 ;
    END
  END b3_r1_b_not
  PIN b3_r0_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 490.870 171.185 492.105 171.565 ;
        RECT 488.845 168.785 492.105 169.165 ;
        RECT 496.275 167.625 509.890 167.925 ;
        RECT 497.470 164.970 501.600 165.270 ;
        RECT 503.975 164.920 508.475 165.230 ;
        RECT 490.730 163.925 494.675 164.260 ;
        RECT 488.825 163.285 492.125 163.665 ;
        RECT 490.640 161.285 492.125 161.665 ;
      LAYER Metal2 ;
        RECT 490.955 161.040 491.270 171.725 ;
        RECT 494.280 163.910 494.660 164.290 ;
        RECT 496.345 163.885 496.655 168.005 ;
        RECT 509.415 167.580 509.710 172.950 ;
      LAYER Metal3 ;
        RECT 509.415 172.495 525.435 172.905 ;
        RECT 494.280 163.900 496.760 164.300 ;
    END
  END b3_r0_b
  PIN b3_r1_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 490.670 151.460 491.905 151.840 ;
        RECT 488.645 149.060 491.905 149.440 ;
        RECT 496.075 147.900 509.690 148.200 ;
        RECT 497.270 145.245 501.400 145.545 ;
        RECT 503.775 145.195 508.275 145.505 ;
        RECT 490.530 144.200 494.475 144.535 ;
        RECT 488.625 143.560 491.925 143.940 ;
        RECT 490.440 141.560 491.925 141.940 ;
      LAYER Metal2 ;
        RECT 490.755 141.315 491.070 152.000 ;
        RECT 494.080 144.185 494.460 144.565 ;
        RECT 496.145 144.160 496.455 148.280 ;
        RECT 509.215 147.855 509.510 153.225 ;
      LAYER Metal3 ;
        RECT 509.215 152.770 525.235 153.180 ;
        RECT 494.080 144.175 496.560 144.575 ;
    END
  END b3_r1_b
  PIN b3_r2_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 471.300 131.715 472.500 132.095 ;
        RECT 471.300 129.415 474.560 129.795 ;
        RECT 471.965 127.500 494.520 127.840 ;
        RECT 495.630 127.510 510.275 127.810 ;
        RECT 471.280 123.915 474.580 124.295 ;
        RECT 498.655 123.835 501.575 124.135 ;
        RECT 505.120 123.820 508.490 124.120 ;
        RECT 471.280 121.915 472.565 122.295 ;
      LAYER Metal2 ;
        RECT 472.125 121.185 472.440 132.235 ;
        RECT 494.100 127.430 494.520 127.890 ;
        RECT 495.600 127.425 496.020 127.885 ;
        RECT 498.690 123.785 498.990 127.845 ;
        RECT 505.180 123.770 505.460 127.860 ;
        RECT 509.945 127.380 510.250 132.855 ;
      LAYER Metal3 ;
        RECT 509.900 132.345 525.380 132.800 ;
        RECT 494.070 127.480 496.095 127.865 ;
    END
  END b3_r2_b_not
  PIN b3_r2_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 490.825 131.815 492.060 132.195 ;
        RECT 488.800 129.415 492.060 129.795 ;
        RECT 496.230 128.255 509.845 128.555 ;
        RECT 497.425 125.600 501.555 125.900 ;
        RECT 503.930 125.550 508.430 125.860 ;
        RECT 490.685 124.555 494.630 124.890 ;
        RECT 488.780 123.915 492.080 124.295 ;
        RECT 490.595 121.915 492.080 122.295 ;
      LAYER Metal2 ;
        RECT 490.910 121.670 491.225 132.355 ;
        RECT 494.235 124.540 494.615 124.920 ;
        RECT 496.300 124.515 496.610 128.635 ;
        RECT 509.370 128.210 509.665 133.580 ;
      LAYER Metal3 ;
        RECT 509.370 133.125 525.390 133.535 ;
        RECT 494.235 124.530 496.715 124.930 ;
    END
  END b3_r2_b
  PIN b3_r3_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 471.300 111.920 472.500 112.300 ;
        RECT 471.300 109.620 474.560 110.000 ;
        RECT 471.965 107.705 494.520 108.045 ;
        RECT 495.630 107.715 510.275 108.015 ;
        RECT 471.280 104.120 474.580 104.500 ;
        RECT 498.655 104.040 501.575 104.340 ;
        RECT 505.120 104.025 508.490 104.325 ;
        RECT 471.280 102.120 472.565 102.500 ;
      LAYER Metal2 ;
        RECT 472.125 101.390 472.440 112.440 ;
        RECT 494.100 107.635 494.520 108.095 ;
        RECT 495.600 107.630 496.020 108.090 ;
        RECT 498.690 103.990 498.990 108.050 ;
        RECT 505.180 103.975 505.460 108.065 ;
        RECT 509.945 107.585 510.250 113.060 ;
      LAYER Metal3 ;
        RECT 509.900 112.550 525.380 113.005 ;
        RECT 494.070 107.685 496.095 108.070 ;
    END
  END b3_r3_b_not
  PIN b3_r3_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 490.825 112.020 492.060 112.400 ;
        RECT 488.800 109.620 492.060 110.000 ;
        RECT 496.230 108.460 509.845 108.760 ;
        RECT 497.425 105.805 501.555 106.105 ;
        RECT 503.930 105.755 508.430 106.065 ;
        RECT 490.685 104.760 494.630 105.095 ;
        RECT 488.780 104.120 492.080 104.500 ;
        RECT 490.595 102.120 492.080 102.500 ;
      LAYER Metal2 ;
        RECT 490.910 101.875 491.225 112.560 ;
        RECT 494.235 104.745 494.615 105.125 ;
        RECT 496.300 104.720 496.610 108.840 ;
        RECT 509.370 108.415 509.665 113.785 ;
      LAYER Metal3 ;
        RECT 509.370 113.330 525.390 113.740 ;
        RECT 494.235 104.735 496.715 105.135 ;
    END
  END b3_r3_b
  PIN b3_r4_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 471.220 92.165 472.420 92.545 ;
        RECT 471.220 89.865 474.480 90.245 ;
        RECT 471.885 87.950 494.440 88.290 ;
        RECT 495.550 87.960 510.195 88.260 ;
        RECT 471.200 84.365 474.500 84.745 ;
        RECT 498.575 84.285 501.495 84.585 ;
        RECT 505.040 84.270 508.410 84.570 ;
        RECT 471.200 82.365 472.485 82.745 ;
      LAYER Metal2 ;
        RECT 472.045 81.635 472.360 92.685 ;
        RECT 494.020 87.880 494.440 88.340 ;
        RECT 495.520 87.875 495.940 88.335 ;
        RECT 498.610 84.235 498.910 88.295 ;
        RECT 505.100 84.220 505.380 88.310 ;
        RECT 509.865 87.830 510.170 93.305 ;
      LAYER Metal3 ;
        RECT 509.820 92.795 525.300 93.250 ;
        RECT 493.990 87.930 496.015 88.315 ;
    END
  END b3_r4_b_not
  PIN b3_r4_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 490.745 92.265 491.980 92.645 ;
        RECT 488.720 89.865 491.980 90.245 ;
        RECT 496.150 88.705 509.765 89.005 ;
        RECT 497.345 86.050 501.475 86.350 ;
        RECT 503.850 86.000 508.350 86.310 ;
        RECT 490.605 85.005 494.550 85.340 ;
        RECT 488.700 84.365 492.000 84.745 ;
        RECT 490.515 82.365 492.000 82.745 ;
      LAYER Metal2 ;
        RECT 490.830 82.120 491.145 92.805 ;
        RECT 494.155 84.990 494.535 85.370 ;
        RECT 496.220 84.965 496.530 89.085 ;
        RECT 509.290 88.660 509.585 94.030 ;
      LAYER Metal3 ;
        RECT 509.290 93.575 525.310 93.985 ;
        RECT 494.155 84.980 496.635 85.380 ;
    END
  END b3_r4_b
  PIN b3_r5_b_not
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 471.325 72.450 472.525 72.830 ;
        RECT 471.325 70.150 474.585 70.530 ;
        RECT 471.990 68.235 494.545 68.575 ;
        RECT 495.655 68.245 510.300 68.545 ;
        RECT 471.305 64.650 474.605 65.030 ;
        RECT 498.680 64.570 501.600 64.870 ;
        RECT 505.145 64.555 508.515 64.855 ;
        RECT 471.305 62.650 472.590 63.030 ;
      LAYER Metal2 ;
        RECT 472.150 61.920 472.465 72.970 ;
        RECT 494.125 68.165 494.545 68.625 ;
        RECT 495.625 68.160 496.045 68.620 ;
        RECT 498.715 64.520 499.015 68.580 ;
        RECT 505.205 64.505 505.485 68.595 ;
        RECT 509.970 68.115 510.275 73.590 ;
      LAYER Metal3 ;
        RECT 509.925 73.080 525.405 73.535 ;
        RECT 494.095 68.215 496.120 68.600 ;
    END
  END b3_r5_b_not
  PIN b3_r5_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 490.850 72.550 492.085 72.930 ;
        RECT 488.825 70.150 492.085 70.530 ;
        RECT 496.255 68.990 509.870 69.290 ;
        RECT 497.450 66.335 501.580 66.635 ;
        RECT 503.955 66.285 508.455 66.595 ;
        RECT 490.710 65.290 494.655 65.625 ;
        RECT 488.805 64.650 492.105 65.030 ;
        RECT 490.620 62.650 492.105 63.030 ;
      LAYER Metal2 ;
        RECT 490.935 62.405 491.250 73.090 ;
        RECT 494.260 65.275 494.640 65.655 ;
        RECT 496.325 65.250 496.635 69.370 ;
        RECT 509.395 68.945 509.690 74.315 ;
      LAYER Metal3 ;
        RECT 509.395 73.860 525.415 74.270 ;
        RECT 494.260 65.265 496.740 65.665 ;
    END
  END b3_r5_b
  PIN p15
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 1257.425 10.840 1257.805 11.220 ;
        RECT 1254.750 10.415 1256.490 10.705 ;
        RECT 1256.105 5.820 1266.510 6.155 ;
        RECT 1256.075 4.500 1257.855 4.790 ;
        RECT 1254.805 3.885 1255.185 4.265 ;
      LAYER Metal2 ;
        RECT 1254.835 3.825 1255.135 10.755 ;
        RECT 1256.145 4.425 1256.445 10.775 ;
        RECT 1257.460 4.455 1257.755 11.280 ;
        RECT 1266.100 5.795 1266.480 6.175 ;
      LAYER Metal3 ;
        RECT 1266.070 5.815 1269.490 6.150 ;
    END
  END p15
  OBS
      LAYER Nwell ;
        RECT -32.455 185.725 -5.800 193.950 ;
      LAYER Pwell ;
        RECT -32.455 178.025 -5.800 185.725 ;
      LAYER Nwell ;
        RECT -82.690 165.990 -56.035 174.215 ;
      LAYER Pwell ;
        RECT -82.690 158.290 -56.035 165.990 ;
      LAYER Nwell ;
        RECT -32.365 166.070 -5.710 174.295 ;
      LAYER Pwell ;
        RECT -32.365 158.370 -5.710 166.070 ;
      LAYER Nwell ;
        RECT 3.385 166.045 62.940 174.270 ;
      LAYER Pwell ;
        RECT 3.385 158.345 34.305 166.045 ;
        RECT 36.285 158.345 62.940 166.045 ;
      LAYER Nwell ;
        RECT 74.875 165.990 132.450 174.215 ;
      LAYER Pwell ;
        RECT 74.875 158.290 132.450 165.990 ;
      LAYER Nwell ;
        RECT 163.805 166.080 190.460 174.305 ;
      LAYER Pwell ;
        RECT 163.805 158.380 190.460 166.080 ;
      LAYER Nwell ;
        RECT 199.750 166.045 259.305 174.270 ;
      LAYER Pwell ;
        RECT 199.750 158.345 230.670 166.045 ;
        RECT 232.650 158.345 259.305 166.045 ;
      LAYER Nwell ;
        RECT 271.240 165.990 328.815 174.215 ;
      LAYER Pwell ;
        RECT 271.240 158.290 328.815 165.990 ;
      LAYER Nwell ;
        RECT 360.195 166.040 386.850 174.265 ;
      LAYER Pwell ;
        RECT 360.195 158.340 386.850 166.040 ;
      LAYER Nwell ;
        RECT 396.150 165.995 455.705 174.220 ;
      LAYER Pwell ;
        RECT 396.150 158.295 427.070 165.995 ;
        RECT 429.050 158.295 455.705 165.995 ;
      LAYER Nwell ;
        RECT 467.640 165.940 525.215 174.165 ;
      LAYER Pwell ;
        RECT 467.640 158.240 525.215 165.940 ;
      LAYER Nwell ;
        RECT 556.515 166.085 583.170 174.310 ;
      LAYER Pwell ;
        RECT 556.515 158.385 583.170 166.085 ;
      LAYER Nwell ;
        RECT 592.525 166.030 652.080 174.255 ;
      LAYER Pwell ;
        RECT 592.525 158.330 623.445 166.030 ;
        RECT 625.425 158.330 652.080 166.030 ;
      LAYER Nwell ;
        RECT 664.015 165.975 721.590 174.200 ;
      LAYER Pwell ;
        RECT 664.015 158.275 721.590 165.975 ;
      LAYER Nwell ;
        RECT 752.880 166.090 779.535 174.315 ;
      LAYER Pwell ;
        RECT 752.880 158.390 779.535 166.090 ;
      LAYER Nwell ;
        RECT 788.865 166.030 848.420 174.255 ;
      LAYER Pwell ;
        RECT 788.865 158.330 819.785 166.030 ;
        RECT 821.765 158.330 848.420 166.030 ;
      LAYER Nwell ;
        RECT 860.355 165.975 917.930 174.200 ;
      LAYER Pwell ;
        RECT 860.355 158.275 917.930 165.975 ;
      LAYER Nwell ;
        RECT 949.265 166.075 975.920 174.300 ;
      LAYER Pwell ;
        RECT 949.265 158.375 975.920 166.075 ;
      LAYER Nwell ;
        RECT 985.205 166.030 1044.760 174.255 ;
      LAYER Pwell ;
        RECT 985.205 158.330 1016.125 166.030 ;
        RECT 1018.105 158.330 1044.760 166.030 ;
      LAYER Nwell ;
        RECT 1056.695 165.975 1114.270 174.200 ;
      LAYER Pwell ;
        RECT 1056.695 158.275 1114.270 165.975 ;
      LAYER Nwell ;
        RECT 1145.590 166.080 1172.245 174.305 ;
      LAYER Pwell ;
        RECT 1145.590 158.380 1172.245 166.080 ;
      LAYER Nwell ;
        RECT 1181.545 166.030 1241.100 174.255 ;
      LAYER Pwell ;
        RECT 1181.545 158.330 1212.465 166.030 ;
        RECT 1214.445 158.330 1241.100 166.030 ;
      LAYER Nwell ;
        RECT 1253.035 165.975 1310.610 174.200 ;
      LAYER Pwell ;
        RECT 1253.035 158.275 1310.610 165.975 ;
      LAYER Nwell ;
        RECT -82.775 146.275 -56.120 154.500 ;
      LAYER Pwell ;
        RECT -82.775 138.575 -56.120 146.275 ;
      LAYER Nwell ;
        RECT -32.450 146.355 -5.795 154.580 ;
      LAYER Pwell ;
        RECT -32.450 138.655 -5.795 146.355 ;
      LAYER Nwell ;
        RECT 3.340 146.355 62.895 154.580 ;
      LAYER Pwell ;
        RECT 3.340 138.655 34.260 146.355 ;
        RECT 36.240 138.655 62.895 146.355 ;
      LAYER Nwell ;
        RECT 74.675 146.265 132.250 154.490 ;
      LAYER Pwell ;
        RECT 74.675 138.565 132.250 146.265 ;
      LAYER Nwell ;
        RECT 163.720 146.365 190.375 154.590 ;
      LAYER Pwell ;
        RECT 163.720 138.665 190.375 146.365 ;
      LAYER Nwell ;
        RECT 199.705 146.355 259.260 154.580 ;
      LAYER Pwell ;
        RECT 199.705 138.655 230.625 146.355 ;
        RECT 232.605 138.655 259.260 146.355 ;
      LAYER Nwell ;
        RECT 271.040 146.265 328.615 154.490 ;
      LAYER Pwell ;
        RECT 271.040 138.565 328.615 146.265 ;
      LAYER Nwell ;
        RECT 360.110 146.325 386.765 154.550 ;
      LAYER Pwell ;
        RECT 360.110 138.625 386.765 146.325 ;
      LAYER Nwell ;
        RECT 396.105 146.305 455.660 154.530 ;
      LAYER Pwell ;
        RECT 396.105 138.605 427.025 146.305 ;
        RECT 429.005 138.605 455.660 146.305 ;
      LAYER Nwell ;
        RECT 467.440 146.215 525.015 154.440 ;
      LAYER Pwell ;
        RECT 467.440 138.515 525.015 146.215 ;
      LAYER Nwell ;
        RECT 556.430 146.370 583.085 154.595 ;
      LAYER Pwell ;
        RECT 556.430 138.670 583.085 146.370 ;
      LAYER Nwell ;
        RECT 592.480 146.340 652.035 154.565 ;
      LAYER Pwell ;
        RECT 592.480 138.640 623.400 146.340 ;
        RECT 625.380 138.640 652.035 146.340 ;
      LAYER Nwell ;
        RECT 663.815 146.250 721.390 154.475 ;
      LAYER Pwell ;
        RECT 663.815 138.550 721.390 146.250 ;
      LAYER Nwell ;
        RECT 752.795 146.375 779.450 154.600 ;
      LAYER Pwell ;
        RECT 752.795 138.675 779.450 146.375 ;
      LAYER Nwell ;
        RECT 788.820 146.340 848.375 154.565 ;
      LAYER Pwell ;
        RECT 788.820 138.640 819.740 146.340 ;
        RECT 821.720 138.640 848.375 146.340 ;
      LAYER Nwell ;
        RECT 860.155 146.250 917.730 154.475 ;
      LAYER Pwell ;
        RECT 860.155 138.550 917.730 146.250 ;
      LAYER Nwell ;
        RECT 949.180 146.360 975.835 154.585 ;
      LAYER Pwell ;
        RECT 949.180 138.660 975.835 146.360 ;
      LAYER Nwell ;
        RECT 985.160 146.340 1044.715 154.565 ;
      LAYER Pwell ;
        RECT 985.160 138.640 1016.080 146.340 ;
        RECT 1018.060 138.640 1044.715 146.340 ;
      LAYER Nwell ;
        RECT 1056.495 146.250 1114.070 154.475 ;
      LAYER Pwell ;
        RECT 1056.495 138.550 1114.070 146.250 ;
      LAYER Nwell ;
        RECT 1145.505 146.365 1172.160 154.590 ;
      LAYER Pwell ;
        RECT 1145.505 138.665 1172.160 146.365 ;
      LAYER Nwell ;
        RECT 1181.500 146.340 1241.055 154.565 ;
      LAYER Pwell ;
        RECT 1181.500 138.640 1212.420 146.340 ;
        RECT 1214.400 138.640 1241.055 146.340 ;
      LAYER Nwell ;
        RECT 1252.835 146.250 1310.410 154.475 ;
      LAYER Pwell ;
        RECT 1252.835 138.550 1310.410 146.250 ;
      LAYER Nwell ;
        RECT -82.715 126.470 -56.060 134.695 ;
      LAYER Pwell ;
        RECT -82.715 118.770 -56.060 126.470 ;
      LAYER Nwell ;
        RECT -32.390 126.550 -5.735 134.775 ;
      LAYER Pwell ;
        RECT -32.390 118.850 -5.735 126.550 ;
      LAYER Nwell ;
        RECT 3.530 126.645 63.085 134.870 ;
      LAYER Pwell ;
        RECT 3.530 118.945 34.450 126.645 ;
        RECT 36.430 118.945 63.085 126.645 ;
      LAYER Nwell ;
        RECT 74.830 126.620 132.405 134.845 ;
      LAYER Pwell ;
        RECT 74.830 118.920 132.405 126.620 ;
      LAYER Nwell ;
        RECT 163.780 126.560 190.435 134.785 ;
      LAYER Pwell ;
        RECT 163.780 118.860 190.435 126.560 ;
      LAYER Nwell ;
        RECT 199.895 126.645 259.450 134.870 ;
      LAYER Pwell ;
        RECT 199.895 118.945 230.815 126.645 ;
        RECT 232.795 118.945 259.450 126.645 ;
      LAYER Nwell ;
        RECT 271.195 126.620 328.770 134.845 ;
      LAYER Pwell ;
        RECT 271.195 118.920 328.770 126.620 ;
      LAYER Nwell ;
        RECT 360.170 126.520 386.825 134.745 ;
      LAYER Pwell ;
        RECT 360.170 118.820 386.825 126.520 ;
      LAYER Nwell ;
        RECT 396.295 126.595 455.850 134.820 ;
      LAYER Pwell ;
        RECT 396.295 118.895 427.215 126.595 ;
        RECT 429.195 118.895 455.850 126.595 ;
      LAYER Nwell ;
        RECT 467.595 126.570 525.170 134.795 ;
      LAYER Pwell ;
        RECT 467.595 118.870 525.170 126.570 ;
      LAYER Nwell ;
        RECT 556.490 126.565 583.145 134.790 ;
      LAYER Pwell ;
        RECT 556.490 118.865 583.145 126.565 ;
      LAYER Nwell ;
        RECT 592.670 126.630 652.225 134.855 ;
      LAYER Pwell ;
        RECT 592.670 118.930 623.590 126.630 ;
        RECT 625.570 118.930 652.225 126.630 ;
      LAYER Nwell ;
        RECT 663.970 126.605 721.545 134.830 ;
      LAYER Pwell ;
        RECT 663.970 118.905 721.545 126.605 ;
      LAYER Nwell ;
        RECT 752.855 126.570 779.510 134.795 ;
      LAYER Pwell ;
        RECT 752.855 118.870 779.510 126.570 ;
      LAYER Nwell ;
        RECT 789.010 126.630 848.565 134.855 ;
      LAYER Pwell ;
        RECT 789.010 118.930 819.930 126.630 ;
        RECT 821.910 118.930 848.565 126.630 ;
      LAYER Nwell ;
        RECT 860.310 126.605 917.885 134.830 ;
      LAYER Pwell ;
        RECT 860.310 118.905 917.885 126.605 ;
      LAYER Nwell ;
        RECT 949.240 126.555 975.895 134.780 ;
      LAYER Pwell ;
        RECT 949.240 118.855 975.895 126.555 ;
      LAYER Nwell ;
        RECT 985.350 126.630 1044.905 134.855 ;
      LAYER Pwell ;
        RECT 985.350 118.930 1016.270 126.630 ;
        RECT 1018.250 118.930 1044.905 126.630 ;
      LAYER Nwell ;
        RECT 1056.650 126.605 1114.225 134.830 ;
      LAYER Pwell ;
        RECT 1056.650 118.905 1114.225 126.605 ;
      LAYER Nwell ;
        RECT 1145.565 126.560 1172.220 134.785 ;
      LAYER Pwell ;
        RECT 1145.565 118.860 1172.220 126.560 ;
      LAYER Nwell ;
        RECT 1181.690 126.630 1241.245 134.855 ;
      LAYER Pwell ;
        RECT 1181.690 118.930 1212.610 126.630 ;
        RECT 1214.590 118.930 1241.245 126.630 ;
      LAYER Nwell ;
        RECT 1252.990 126.605 1310.565 134.830 ;
      LAYER Pwell ;
        RECT 1252.990 118.905 1310.565 126.605 ;
      LAYER Nwell ;
        RECT -82.785 106.700 -56.130 114.925 ;
      LAYER Pwell ;
        RECT -82.785 99.000 -56.130 106.700 ;
      LAYER Nwell ;
        RECT -32.460 106.780 -5.805 115.005 ;
      LAYER Pwell ;
        RECT -32.460 99.080 -5.805 106.780 ;
      LAYER Nwell ;
        RECT 3.335 106.805 62.890 115.030 ;
      LAYER Pwell ;
        RECT 3.335 99.105 34.255 106.805 ;
        RECT 36.235 99.105 62.890 106.805 ;
      LAYER Nwell ;
        RECT 74.830 106.825 132.405 115.050 ;
      LAYER Pwell ;
        RECT 74.830 99.125 132.405 106.825 ;
      LAYER Nwell ;
        RECT 163.710 106.790 190.365 115.015 ;
      LAYER Pwell ;
        RECT 163.710 99.090 190.365 106.790 ;
      LAYER Nwell ;
        RECT 199.700 106.805 259.255 115.030 ;
      LAYER Pwell ;
        RECT 199.700 99.105 230.620 106.805 ;
        RECT 232.600 99.105 259.255 106.805 ;
      LAYER Nwell ;
        RECT 271.195 106.825 328.770 115.050 ;
      LAYER Pwell ;
        RECT 271.195 99.125 328.770 106.825 ;
      LAYER Nwell ;
        RECT 360.100 106.750 386.755 114.975 ;
      LAYER Pwell ;
        RECT 360.100 99.050 386.755 106.750 ;
      LAYER Nwell ;
        RECT 396.100 106.755 455.655 114.980 ;
      LAYER Pwell ;
        RECT 396.100 99.055 427.020 106.755 ;
        RECT 429.000 99.055 455.655 106.755 ;
      LAYER Nwell ;
        RECT 467.595 106.775 525.170 115.000 ;
      LAYER Pwell ;
        RECT 467.595 99.075 525.170 106.775 ;
      LAYER Nwell ;
        RECT 556.420 106.795 583.075 115.020 ;
      LAYER Pwell ;
        RECT 556.420 99.095 583.075 106.795 ;
      LAYER Nwell ;
        RECT 592.475 106.790 652.030 115.015 ;
      LAYER Pwell ;
        RECT 592.475 99.090 623.395 106.790 ;
        RECT 625.375 99.090 652.030 106.790 ;
      LAYER Nwell ;
        RECT 663.970 106.810 721.545 115.035 ;
      LAYER Pwell ;
        RECT 663.970 99.110 721.545 106.810 ;
      LAYER Nwell ;
        RECT 752.785 106.800 779.440 115.025 ;
      LAYER Pwell ;
        RECT 752.785 99.100 779.440 106.800 ;
      LAYER Nwell ;
        RECT 788.815 106.790 848.370 115.015 ;
      LAYER Pwell ;
        RECT 788.815 99.090 819.735 106.790 ;
        RECT 821.715 99.090 848.370 106.790 ;
      LAYER Nwell ;
        RECT 860.310 106.810 917.885 115.035 ;
      LAYER Pwell ;
        RECT 860.310 99.110 917.885 106.810 ;
      LAYER Nwell ;
        RECT 949.170 106.785 975.825 115.010 ;
      LAYER Pwell ;
        RECT 949.170 99.085 975.825 106.785 ;
      LAYER Nwell ;
        RECT 985.155 106.790 1044.710 115.015 ;
      LAYER Pwell ;
        RECT 985.155 99.090 1016.075 106.790 ;
        RECT 1018.055 99.090 1044.710 106.790 ;
      LAYER Nwell ;
        RECT 1056.650 106.810 1114.225 115.035 ;
      LAYER Pwell ;
        RECT 1056.650 99.110 1114.225 106.810 ;
      LAYER Nwell ;
        RECT 1145.495 106.790 1172.150 115.015 ;
      LAYER Pwell ;
        RECT 1145.495 99.090 1172.150 106.790 ;
      LAYER Nwell ;
        RECT 1181.495 106.790 1241.050 115.015 ;
      LAYER Pwell ;
        RECT 1181.495 99.090 1212.415 106.790 ;
        RECT 1214.395 99.090 1241.050 106.790 ;
      LAYER Nwell ;
        RECT 1252.990 106.810 1310.565 115.035 ;
      LAYER Pwell ;
        RECT 1252.990 99.110 1310.565 106.810 ;
      LAYER Nwell ;
        RECT -82.755 86.975 -56.100 95.200 ;
      LAYER Pwell ;
        RECT -82.755 79.275 -56.100 86.975 ;
      LAYER Nwell ;
        RECT -32.430 87.055 -5.775 95.280 ;
      LAYER Pwell ;
        RECT -32.430 79.355 -5.775 87.055 ;
      LAYER Nwell ;
        RECT 3.205 87.095 62.760 95.320 ;
      LAYER Pwell ;
        RECT 3.205 79.395 34.125 87.095 ;
        RECT 36.105 79.395 62.760 87.095 ;
      LAYER Nwell ;
        RECT 74.750 87.070 132.325 95.295 ;
      LAYER Pwell ;
        RECT 74.750 79.370 132.325 87.070 ;
      LAYER Nwell ;
        RECT 163.740 87.065 190.395 95.290 ;
      LAYER Pwell ;
        RECT 163.740 79.365 190.395 87.065 ;
      LAYER Nwell ;
        RECT 199.570 87.095 259.125 95.320 ;
      LAYER Pwell ;
        RECT 199.570 79.395 230.490 87.095 ;
        RECT 232.470 79.395 259.125 87.095 ;
      LAYER Nwell ;
        RECT 271.115 87.070 328.690 95.295 ;
      LAYER Pwell ;
        RECT 271.115 79.370 328.690 87.070 ;
      LAYER Nwell ;
        RECT 360.130 87.025 386.785 95.250 ;
      LAYER Pwell ;
        RECT 360.130 79.325 386.785 87.025 ;
      LAYER Nwell ;
        RECT 395.970 87.045 455.525 95.270 ;
      LAYER Pwell ;
        RECT 395.970 79.345 426.890 87.045 ;
        RECT 428.870 79.345 455.525 87.045 ;
      LAYER Nwell ;
        RECT 467.515 87.020 525.090 95.245 ;
      LAYER Pwell ;
        RECT 467.515 79.320 525.090 87.020 ;
      LAYER Nwell ;
        RECT 556.450 87.070 583.105 95.295 ;
      LAYER Pwell ;
        RECT 556.450 79.370 583.105 87.070 ;
      LAYER Nwell ;
        RECT 592.345 87.080 651.900 95.305 ;
      LAYER Pwell ;
        RECT 592.345 79.380 623.265 87.080 ;
        RECT 625.245 79.380 651.900 87.080 ;
      LAYER Nwell ;
        RECT 663.890 87.055 721.465 95.280 ;
      LAYER Pwell ;
        RECT 663.890 79.355 721.465 87.055 ;
      LAYER Nwell ;
        RECT 752.815 87.075 779.470 95.300 ;
      LAYER Pwell ;
        RECT 752.815 79.375 779.470 87.075 ;
      LAYER Nwell ;
        RECT 788.685 87.080 848.240 95.305 ;
      LAYER Pwell ;
        RECT 788.685 79.380 819.605 87.080 ;
        RECT 821.585 79.380 848.240 87.080 ;
      LAYER Nwell ;
        RECT 860.230 87.055 917.805 95.280 ;
      LAYER Pwell ;
        RECT 860.230 79.355 917.805 87.055 ;
      LAYER Nwell ;
        RECT 949.200 87.060 975.855 95.285 ;
      LAYER Pwell ;
        RECT 949.200 79.360 975.855 87.060 ;
      LAYER Nwell ;
        RECT 985.025 87.080 1044.580 95.305 ;
      LAYER Pwell ;
        RECT 985.025 79.380 1015.945 87.080 ;
        RECT 1017.925 79.380 1044.580 87.080 ;
      LAYER Nwell ;
        RECT 1056.570 87.055 1114.145 95.280 ;
      LAYER Pwell ;
        RECT 1056.570 79.355 1114.145 87.055 ;
      LAYER Nwell ;
        RECT 1145.525 87.065 1172.180 95.290 ;
      LAYER Pwell ;
        RECT 1145.525 79.365 1172.180 87.065 ;
      LAYER Nwell ;
        RECT 1181.365 87.080 1240.920 95.305 ;
      LAYER Pwell ;
        RECT 1181.365 79.380 1212.285 87.080 ;
        RECT 1214.265 79.380 1240.920 87.080 ;
      LAYER Nwell ;
        RECT 1252.910 87.055 1310.485 95.280 ;
      LAYER Pwell ;
        RECT 1252.910 79.355 1310.485 87.055 ;
      LAYER Nwell ;
        RECT -82.825 67.145 -56.170 75.370 ;
      LAYER Pwell ;
        RECT -82.825 59.445 -56.170 67.145 ;
      LAYER Nwell ;
        RECT -32.500 67.225 -5.845 75.450 ;
      LAYER Pwell ;
        RECT -32.500 59.525 -5.845 67.225 ;
      LAYER Nwell ;
        RECT 3.335 67.335 62.890 75.560 ;
      LAYER Pwell ;
        RECT 3.335 59.635 34.255 67.335 ;
        RECT 36.235 59.635 62.890 67.335 ;
      LAYER Nwell ;
        RECT 74.855 67.355 132.430 75.580 ;
      LAYER Pwell ;
        RECT 74.855 59.655 132.430 67.355 ;
      LAYER Nwell ;
        RECT 163.670 67.235 190.325 75.460 ;
      LAYER Pwell ;
        RECT 163.670 59.535 190.325 67.235 ;
      LAYER Nwell ;
        RECT 199.700 67.335 259.255 75.560 ;
      LAYER Pwell ;
        RECT 199.700 59.635 230.620 67.335 ;
        RECT 232.600 59.635 259.255 67.335 ;
      LAYER Nwell ;
        RECT 271.220 67.355 328.795 75.580 ;
      LAYER Pwell ;
        RECT 271.220 59.655 328.795 67.355 ;
      LAYER Nwell ;
        RECT 360.060 67.195 386.715 75.420 ;
      LAYER Pwell ;
        RECT 360.060 59.495 386.715 67.195 ;
      LAYER Nwell ;
        RECT 396.100 67.285 455.655 75.510 ;
      LAYER Pwell ;
        RECT 396.100 59.585 427.020 67.285 ;
        RECT 429.000 59.585 455.655 67.285 ;
      LAYER Nwell ;
        RECT 467.620 67.305 525.195 75.530 ;
      LAYER Pwell ;
        RECT 467.620 59.605 525.195 67.305 ;
      LAYER Nwell ;
        RECT 556.380 67.240 583.035 75.465 ;
      LAYER Pwell ;
        RECT 556.380 59.540 583.035 67.240 ;
      LAYER Nwell ;
        RECT 592.475 67.320 652.030 75.545 ;
      LAYER Pwell ;
        RECT 592.475 59.620 623.395 67.320 ;
        RECT 625.375 59.620 652.030 67.320 ;
      LAYER Nwell ;
        RECT 663.995 67.340 721.570 75.565 ;
      LAYER Pwell ;
        RECT 663.995 59.640 721.570 67.340 ;
      LAYER Nwell ;
        RECT 752.745 67.245 779.400 75.470 ;
      LAYER Pwell ;
        RECT 752.745 59.545 779.400 67.245 ;
      LAYER Nwell ;
        RECT 788.815 67.320 848.370 75.545 ;
      LAYER Pwell ;
        RECT 788.815 59.620 819.735 67.320 ;
        RECT 821.715 59.620 848.370 67.320 ;
      LAYER Nwell ;
        RECT 860.335 67.340 917.910 75.565 ;
      LAYER Pwell ;
        RECT 860.335 59.640 917.910 67.340 ;
      LAYER Nwell ;
        RECT 949.130 67.230 975.785 75.455 ;
      LAYER Pwell ;
        RECT 949.130 59.530 975.785 67.230 ;
      LAYER Nwell ;
        RECT 985.155 67.320 1044.710 75.545 ;
      LAYER Pwell ;
        RECT 985.155 59.620 1016.075 67.320 ;
        RECT 1018.055 59.620 1044.710 67.320 ;
      LAYER Nwell ;
        RECT 1056.675 67.340 1114.250 75.565 ;
      LAYER Pwell ;
        RECT 1056.675 59.640 1114.250 67.340 ;
      LAYER Nwell ;
        RECT 1145.455 67.235 1172.110 75.460 ;
      LAYER Pwell ;
        RECT 1145.455 59.535 1172.110 67.235 ;
      LAYER Nwell ;
        RECT 1181.495 67.320 1241.050 75.545 ;
      LAYER Pwell ;
        RECT 1181.495 59.620 1212.415 67.320 ;
        RECT 1214.395 59.620 1241.050 67.320 ;
      LAYER Nwell ;
        RECT 1253.015 67.340 1310.590 75.565 ;
      LAYER Pwell ;
        RECT 1253.015 59.640 1310.590 67.340 ;
      LAYER Nwell ;
        RECT -82.755 47.425 -56.100 55.650 ;
      LAYER Pwell ;
        RECT -82.755 39.725 -56.100 47.425 ;
      LAYER Nwell ;
        RECT -32.430 47.505 -5.775 55.730 ;
      LAYER Pwell ;
        RECT -32.430 39.805 -5.775 47.505 ;
      LAYER Nwell ;
        RECT 3.285 47.525 62.840 55.750 ;
      LAYER Pwell ;
        RECT 3.285 39.825 34.205 47.525 ;
        RECT 36.185 39.825 62.840 47.525 ;
      LAYER Nwell ;
        RECT 74.855 47.385 132.430 55.610 ;
      LAYER Pwell ;
        RECT 74.855 39.685 132.430 47.385 ;
      LAYER Nwell ;
        RECT 163.740 47.515 190.395 55.740 ;
      LAYER Pwell ;
        RECT 163.740 39.815 190.395 47.515 ;
      LAYER Nwell ;
        RECT 199.650 47.525 259.205 55.750 ;
      LAYER Pwell ;
        RECT 199.650 39.825 230.570 47.525 ;
        RECT 232.550 39.825 259.205 47.525 ;
      LAYER Nwell ;
        RECT 271.220 47.385 328.795 55.610 ;
      LAYER Pwell ;
        RECT 271.220 39.685 328.795 47.385 ;
      LAYER Nwell ;
        RECT 360.130 47.475 386.785 55.700 ;
      LAYER Pwell ;
        RECT 360.130 39.775 386.785 47.475 ;
      LAYER Nwell ;
        RECT 396.050 47.475 455.605 55.700 ;
      LAYER Pwell ;
        RECT 396.050 39.775 426.970 47.475 ;
        RECT 428.950 39.775 455.605 47.475 ;
      LAYER Nwell ;
        RECT 467.620 47.335 525.195 55.560 ;
      LAYER Pwell ;
        RECT 467.620 39.635 525.195 47.335 ;
      LAYER Nwell ;
        RECT 556.450 47.520 583.105 55.745 ;
      LAYER Pwell ;
        RECT 556.450 39.820 583.105 47.520 ;
      LAYER Nwell ;
        RECT 592.425 47.510 651.980 55.735 ;
      LAYER Pwell ;
        RECT 592.425 39.810 623.345 47.510 ;
        RECT 625.325 39.810 651.980 47.510 ;
      LAYER Nwell ;
        RECT 663.995 47.370 721.570 55.595 ;
      LAYER Pwell ;
        RECT 663.995 39.670 721.570 47.370 ;
      LAYER Nwell ;
        RECT 752.815 47.525 779.470 55.750 ;
      LAYER Pwell ;
        RECT 752.815 39.825 779.470 47.525 ;
      LAYER Nwell ;
        RECT 788.765 47.510 848.320 55.735 ;
      LAYER Pwell ;
        RECT 788.765 39.810 819.685 47.510 ;
        RECT 821.665 39.810 848.320 47.510 ;
      LAYER Nwell ;
        RECT 860.335 47.370 917.910 55.595 ;
      LAYER Pwell ;
        RECT 860.335 39.670 917.910 47.370 ;
      LAYER Nwell ;
        RECT 949.200 47.510 975.855 55.735 ;
      LAYER Pwell ;
        RECT 949.200 39.810 975.855 47.510 ;
      LAYER Nwell ;
        RECT 985.105 47.510 1044.660 55.735 ;
      LAYER Pwell ;
        RECT 985.105 39.810 1016.025 47.510 ;
        RECT 1018.005 39.810 1044.660 47.510 ;
      LAYER Nwell ;
        RECT 1056.675 47.370 1114.250 55.595 ;
      LAYER Pwell ;
        RECT 1056.675 39.670 1114.250 47.370 ;
      LAYER Nwell ;
        RECT 1145.525 47.515 1172.180 55.740 ;
      LAYER Pwell ;
        RECT 1145.525 39.815 1172.180 47.515 ;
      LAYER Nwell ;
        RECT 1181.445 47.510 1241.000 55.735 ;
      LAYER Pwell ;
        RECT 1181.445 39.810 1212.365 47.510 ;
        RECT 1214.345 39.810 1241.000 47.510 ;
      LAYER Nwell ;
        RECT 1253.015 47.370 1310.590 55.595 ;
      LAYER Pwell ;
        RECT 1253.015 39.670 1310.590 47.370 ;
      LAYER Nwell ;
        RECT -82.750 27.615 -56.095 35.840 ;
      LAYER Pwell ;
        RECT -82.750 19.915 -56.095 27.615 ;
      LAYER Nwell ;
        RECT 3.255 27.730 62.810 35.955 ;
      LAYER Pwell ;
        RECT 3.255 20.030 34.175 27.730 ;
        RECT 36.155 20.030 62.810 27.730 ;
      LAYER Nwell ;
        RECT 74.855 27.720 132.430 35.945 ;
      LAYER Pwell ;
        RECT 74.855 20.020 132.430 27.720 ;
      LAYER Nwell ;
        RECT 163.715 27.785 190.370 36.010 ;
      LAYER Pwell ;
        RECT 163.715 20.085 190.370 27.785 ;
      LAYER Nwell ;
        RECT 199.620 27.730 259.175 35.955 ;
      LAYER Pwell ;
        RECT 199.620 20.030 230.540 27.730 ;
        RECT 232.520 20.030 259.175 27.730 ;
      LAYER Nwell ;
        RECT 271.220 27.720 328.795 35.945 ;
      LAYER Pwell ;
        RECT 271.220 20.020 328.795 27.720 ;
      LAYER Nwell ;
        RECT 360.105 27.745 386.760 35.970 ;
      LAYER Pwell ;
        RECT 360.105 20.045 386.760 27.745 ;
      LAYER Nwell ;
        RECT 396.020 27.680 455.575 35.905 ;
      LAYER Pwell ;
        RECT 396.020 19.980 426.940 27.680 ;
        RECT 428.920 19.980 455.575 27.680 ;
      LAYER Nwell ;
        RECT 467.620 27.670 525.195 35.895 ;
      LAYER Pwell ;
        RECT 467.620 19.970 525.195 27.670 ;
      LAYER Nwell ;
        RECT 556.425 27.790 583.080 36.015 ;
      LAYER Pwell ;
        RECT 556.425 20.090 583.080 27.790 ;
      LAYER Nwell ;
        RECT 592.395 27.715 651.950 35.940 ;
      LAYER Pwell ;
        RECT 592.395 20.015 623.315 27.715 ;
        RECT 625.295 20.015 651.950 27.715 ;
      LAYER Nwell ;
        RECT 663.995 27.705 721.570 35.930 ;
      LAYER Pwell ;
        RECT 663.995 20.005 721.570 27.705 ;
      LAYER Nwell ;
        RECT 752.790 27.795 779.445 36.020 ;
      LAYER Pwell ;
        RECT 752.790 20.095 779.445 27.795 ;
      LAYER Nwell ;
        RECT 788.735 27.715 848.290 35.940 ;
      LAYER Pwell ;
        RECT 788.735 20.015 819.655 27.715 ;
        RECT 821.635 20.015 848.290 27.715 ;
      LAYER Nwell ;
        RECT 860.335 27.705 917.910 35.930 ;
      LAYER Pwell ;
        RECT 860.335 20.005 917.910 27.705 ;
      LAYER Nwell ;
        RECT 949.175 27.780 975.830 36.005 ;
      LAYER Pwell ;
        RECT 949.175 20.080 975.830 27.780 ;
      LAYER Nwell ;
        RECT 985.075 27.715 1044.630 35.940 ;
      LAYER Pwell ;
        RECT 985.075 20.015 1015.995 27.715 ;
        RECT 1017.975 20.015 1044.630 27.715 ;
      LAYER Nwell ;
        RECT 1056.675 27.705 1114.250 35.930 ;
      LAYER Pwell ;
        RECT 1056.675 20.005 1114.250 27.705 ;
      LAYER Nwell ;
        RECT 1145.500 27.785 1172.155 36.010 ;
      LAYER Pwell ;
        RECT 1145.500 20.085 1172.155 27.785 ;
      LAYER Nwell ;
        RECT 1181.415 27.715 1240.970 35.940 ;
      LAYER Pwell ;
        RECT 1181.415 20.015 1212.335 27.715 ;
        RECT 1214.315 20.015 1240.970 27.715 ;
      LAYER Nwell ;
        RECT 1253.015 27.705 1310.590 35.930 ;
      LAYER Pwell ;
        RECT 1253.015 20.005 1310.590 27.705 ;
      LAYER Metal1 ;
        RECT -31.235 193.050 -5.800 193.950 ;
        RECT -25.795 190.655 -23.520 191.165 ;
        RECT -20.895 190.655 -18.595 191.165 ;
        RECT -16.300 190.655 -14.020 191.165 ;
        RECT -24.750 188.570 -21.490 188.950 ;
        RECT -15.250 188.570 -11.990 188.950 ;
        RECT -24.770 183.070 -21.470 183.450 ;
        RECT -15.270 183.070 -11.970 183.450 ;
        RECT -27.265 180.390 -25.745 180.750 ;
        RECT -32.455 178.025 -5.800 178.925 ;
        RECT -81.470 173.315 -56.035 174.215 ;
        RECT -31.145 173.395 -5.710 174.295 ;
        RECT 3.815 174.215 76.205 174.270 ;
        RECT 3.815 173.370 132.450 174.215 ;
        RECT 165.025 173.405 190.460 174.305 ;
        RECT 200.180 174.215 272.570 174.270 ;
        RECT 200.180 173.370 328.815 174.215 ;
        RECT -78.985 171.135 -77.785 171.515 ;
        RECT -76.030 170.920 -73.755 171.430 ;
        RECT -71.130 170.920 -68.830 171.430 ;
        RECT -66.535 170.920 -64.255 171.430 ;
        RECT -59.460 171.235 -58.225 171.615 ;
        RECT -28.660 171.215 -27.460 171.595 ;
        RECT -25.705 171.000 -23.430 171.510 ;
        RECT -20.805 171.000 -18.505 171.510 ;
        RECT -16.210 171.000 -13.930 171.510 ;
        RECT -9.135 171.315 -7.900 171.695 ;
        RECT -78.985 168.835 -75.725 169.215 ;
        RECT -74.985 168.835 -71.725 169.215 ;
        RECT -65.485 168.835 -62.225 169.215 ;
        RECT -61.485 168.835 -58.225 169.215 ;
        RECT -28.660 168.915 -25.400 169.295 ;
        RECT -24.660 168.915 -21.400 169.295 ;
        RECT -15.160 168.915 -11.900 169.295 ;
        RECT -11.160 168.915 -7.900 169.295 ;
        RECT -78.320 167.250 -56.035 167.260 ;
        RECT -78.320 166.920 -54.495 167.250 ;
        RECT -27.995 167.000 -1.700 167.340 ;
        RECT -56.255 166.900 -54.495 166.920 ;
        RECT 4.185 166.210 4.565 173.370 ;
        RECT 6.015 169.155 9.390 169.555 ;
        RECT 9.760 168.915 10.140 169.295 ;
        RECT 12.475 168.955 12.855 169.335 ;
        RECT 16.660 168.905 17.040 169.285 ;
        RECT 7.085 168.490 8.825 168.780 ;
        RECT 10.875 168.440 12.075 168.730 ;
        RECT 13.585 168.410 16.195 168.835 ;
        RECT 17.795 168.505 18.175 168.885 ;
        RECT 5.330 167.730 18.895 168.045 ;
        RECT 5.325 166.985 18.885 167.285 ;
        RECT 5.345 166.270 12.070 166.570 ;
        RECT 15.770 165.970 18.875 166.245 ;
        RECT 19.645 166.210 20.025 173.370 ;
        RECT 76.095 173.315 132.450 173.370 ;
        RECT 36.285 172.330 73.835 172.385 ;
        RECT 36.285 172.100 101.855 172.330 ;
        RECT 73.080 172.045 101.855 172.100 ;
        RECT 103.525 172.025 110.230 172.325 ;
        RECT 37.795 171.190 39.250 171.570 ;
        RECT 39.990 171.190 41.190 171.570 ;
        RECT 42.945 170.975 45.220 171.485 ;
        RECT 47.845 170.975 50.145 171.485 ;
        RECT 52.440 170.975 54.720 171.485 ;
        RECT 59.515 171.290 60.750 171.670 ;
        RECT 61.490 171.290 62.770 171.670 ;
        RECT 76.385 171.135 77.840 171.515 ;
        RECT 60.930 170.935 61.310 170.970 ;
        RECT 39.430 170.830 39.810 170.870 ;
        RECT 39.360 170.525 42.195 170.830 ;
        RECT 58.175 170.625 61.310 170.935 ;
        RECT 81.535 170.920 83.810 171.430 ;
        RECT 86.435 170.920 88.735 171.430 ;
        RECT 91.030 170.920 93.310 171.430 ;
        RECT 100.080 171.235 101.360 171.615 ;
        RECT 99.520 170.880 99.900 170.915 ;
        RECT 78.020 170.775 78.400 170.815 ;
        RECT 60.930 170.590 61.310 170.625 ;
        RECT 39.430 170.490 39.810 170.525 ;
        RECT 77.950 170.470 80.785 170.775 ;
        RECT 96.765 170.570 99.900 170.880 ;
        RECT 99.520 170.535 99.900 170.570 ;
        RECT 78.020 170.435 78.400 170.470 ;
        RECT 25.220 168.915 25.600 169.295 ;
        RECT 32.120 168.905 32.500 169.285 ;
        RECT 37.955 168.890 39.250 169.270 ;
        RECT 39.990 168.890 43.250 169.270 ;
        RECT 43.990 168.890 47.250 169.270 ;
        RECT 47.990 168.890 49.175 169.270 ;
        RECT 51.440 168.890 52.750 169.270 ;
        RECT 53.490 168.890 56.750 169.270 ;
        RECT 57.490 168.890 60.750 169.270 ;
        RECT 61.490 168.890 62.505 169.270 ;
        RECT 76.545 168.835 77.840 169.215 ;
        RECT 82.580 168.835 85.840 169.215 ;
        RECT 86.580 168.835 87.765 169.215 ;
        RECT 90.030 168.835 91.340 169.215 ;
        RECT 92.080 168.835 95.340 169.215 ;
        RECT 100.080 168.835 101.095 169.215 ;
        RECT 104.160 169.080 107.575 169.500 ;
        RECT 110.620 168.900 111.000 169.280 ;
        RECT 22.545 168.490 24.285 168.780 ;
        RECT 29.045 168.410 31.640 168.785 ;
        RECT 39.430 168.190 39.810 168.570 ;
        RECT 43.430 168.190 43.810 168.570 ;
        RECT 47.430 168.525 47.810 168.570 ;
        RECT 52.930 168.525 53.310 168.570 ;
        RECT 47.380 168.210 53.315 168.525 ;
        RECT 47.430 168.190 47.810 168.210 ;
        RECT 52.930 168.190 53.310 168.210 ;
        RECT 56.930 168.190 57.310 168.570 ;
        RECT 60.930 168.190 61.310 168.570 ;
        RECT 78.020 168.135 78.400 168.515 ;
        RECT 82.020 168.135 82.400 168.515 ;
        RECT 86.020 168.470 86.400 168.515 ;
        RECT 91.520 168.470 91.900 168.515 ;
        RECT 85.970 168.155 91.905 168.470 ;
        RECT 86.020 168.135 86.400 168.155 ;
        RECT 91.520 168.135 91.900 168.155 ;
        RECT 95.520 168.135 95.900 168.515 ;
        RECT 99.520 168.135 99.900 168.515 ;
        RECT 109.020 168.385 110.220 168.675 ;
        RECT 115.940 168.450 116.320 168.830 ;
        RECT 20.785 167.730 34.610 168.030 ;
        RECT 36.285 167.565 52.295 167.940 ;
        RECT 70.110 167.510 90.885 167.885 ;
        RECT 20.790 166.985 39.210 167.285 ;
        RECT 40.655 166.975 67.965 167.315 ;
        RECT 31.230 165.970 34.980 166.245 ;
        RECT 36.285 166.210 62.515 166.600 ;
        RECT 69.140 166.155 101.105 166.545 ;
        RECT 117.790 166.155 118.170 173.315 ;
        RECT 167.510 171.225 168.710 171.605 ;
        RECT 119.030 170.855 125.770 171.155 ;
        RECT 170.465 171.010 172.740 171.520 ;
        RECT 175.365 171.010 177.665 171.520 ;
        RECT 179.960 171.010 182.240 171.520 ;
        RECT 187.035 171.325 188.270 171.705 ;
        RECT 119.620 169.060 123.075 169.500 ;
        RECT 126.080 168.900 126.460 169.280 ;
        RECT 167.510 168.925 170.770 169.305 ;
        RECT 171.510 168.925 174.770 169.305 ;
        RECT 181.010 168.925 184.270 169.305 ;
        RECT 185.010 168.925 188.270 169.305 ;
        RECT 124.480 168.385 125.680 168.675 ;
        RECT 131.400 168.450 131.780 168.830 ;
        RECT 168.175 167.010 194.470 167.350 ;
        RECT 200.550 166.210 200.930 173.370 ;
        RECT 202.380 169.155 205.755 169.555 ;
        RECT 206.125 168.915 206.505 169.295 ;
        RECT 208.840 168.955 209.220 169.335 ;
        RECT 213.025 168.905 213.405 169.285 ;
        RECT 203.450 168.490 205.190 168.780 ;
        RECT 207.240 168.440 208.440 168.730 ;
        RECT 209.950 168.410 212.560 168.835 ;
        RECT 214.160 168.505 214.540 168.885 ;
        RECT 201.695 167.730 215.260 168.045 ;
        RECT 201.690 166.985 215.250 167.285 ;
        RECT 201.710 166.270 208.435 166.570 ;
        RECT 212.135 165.970 215.240 166.245 ;
        RECT 216.010 166.210 216.390 173.370 ;
        RECT 272.460 173.315 328.815 173.370 ;
        RECT 361.415 173.365 386.850 174.265 ;
        RECT 396.580 174.165 468.970 174.220 ;
        RECT 396.580 173.320 525.215 174.165 ;
        RECT 557.735 173.410 583.170 174.310 ;
        RECT 592.955 174.200 665.345 174.255 ;
        RECT 592.955 173.355 721.590 174.200 ;
        RECT 754.100 173.415 779.535 174.315 ;
        RECT 789.295 174.200 861.685 174.255 ;
        RECT 789.295 173.355 917.930 174.200 ;
        RECT 950.485 173.400 975.920 174.300 ;
        RECT 985.635 174.200 1058.025 174.255 ;
        RECT 985.635 173.355 1114.270 174.200 ;
        RECT 1146.810 173.405 1172.245 174.305 ;
        RECT 1181.975 174.200 1254.365 174.255 ;
        RECT 1181.975 173.355 1310.610 174.200 ;
        RECT 232.650 172.330 270.200 172.385 ;
        RECT 232.650 172.100 298.220 172.330 ;
        RECT 269.445 172.045 298.220 172.100 ;
        RECT 299.890 172.025 306.595 172.325 ;
        RECT 234.160 171.190 235.615 171.570 ;
        RECT 236.355 171.190 237.555 171.570 ;
        RECT 239.310 170.975 241.585 171.485 ;
        RECT 244.210 170.975 246.510 171.485 ;
        RECT 248.805 170.975 251.085 171.485 ;
        RECT 255.880 171.290 257.115 171.670 ;
        RECT 257.855 171.290 259.135 171.670 ;
        RECT 272.750 171.135 274.205 171.515 ;
        RECT 257.295 170.935 257.675 170.970 ;
        RECT 235.795 170.830 236.175 170.870 ;
        RECT 235.725 170.525 238.560 170.830 ;
        RECT 254.540 170.625 257.675 170.935 ;
        RECT 277.900 170.920 280.175 171.430 ;
        RECT 282.800 170.920 285.100 171.430 ;
        RECT 287.395 170.920 289.675 171.430 ;
        RECT 296.445 171.235 297.725 171.615 ;
        RECT 295.885 170.880 296.265 170.915 ;
        RECT 274.385 170.775 274.765 170.815 ;
        RECT 257.295 170.590 257.675 170.625 ;
        RECT 235.795 170.490 236.175 170.525 ;
        RECT 274.315 170.470 277.150 170.775 ;
        RECT 293.130 170.570 296.265 170.880 ;
        RECT 295.885 170.535 296.265 170.570 ;
        RECT 274.385 170.435 274.765 170.470 ;
        RECT 217.840 169.115 221.245 169.555 ;
        RECT 221.585 168.915 221.965 169.295 ;
        RECT 224.300 168.955 224.680 169.335 ;
        RECT 228.485 168.905 228.865 169.285 ;
        RECT 234.320 168.890 235.615 169.270 ;
        RECT 236.355 168.890 239.615 169.270 ;
        RECT 240.355 168.890 243.615 169.270 ;
        RECT 244.355 168.890 245.540 169.270 ;
        RECT 247.805 168.890 249.115 169.270 ;
        RECT 249.855 168.890 253.115 169.270 ;
        RECT 253.855 168.890 257.115 169.270 ;
        RECT 257.855 168.890 258.870 169.270 ;
        RECT 218.910 168.490 220.650 168.780 ;
        RECT 222.700 168.440 223.900 168.730 ;
        RECT 225.410 168.410 228.005 168.785 ;
        RECT 229.620 168.505 230.000 168.885 ;
        RECT 272.910 168.835 274.205 169.215 ;
        RECT 278.945 168.835 282.205 169.215 ;
        RECT 282.945 168.835 284.130 169.215 ;
        RECT 286.395 168.835 287.705 169.215 ;
        RECT 288.445 168.835 291.705 169.215 ;
        RECT 296.445 168.835 297.460 169.215 ;
        RECT 300.525 169.080 303.940 169.500 ;
        RECT 304.270 168.860 304.650 169.240 ;
        RECT 306.985 168.900 307.365 169.280 ;
        RECT 311.170 168.850 311.550 169.230 ;
        RECT 235.795 168.190 236.175 168.570 ;
        RECT 239.795 168.190 240.175 168.570 ;
        RECT 243.795 168.525 244.175 168.570 ;
        RECT 249.295 168.525 249.675 168.570 ;
        RECT 243.745 168.210 249.680 168.525 ;
        RECT 243.795 168.190 244.175 168.210 ;
        RECT 249.295 168.190 249.675 168.210 ;
        RECT 253.295 168.190 253.675 168.570 ;
        RECT 257.295 168.190 257.675 168.570 ;
        RECT 274.385 168.135 274.765 168.515 ;
        RECT 278.385 168.135 278.765 168.515 ;
        RECT 282.385 168.470 282.765 168.515 ;
        RECT 287.885 168.470 288.265 168.515 ;
        RECT 282.335 168.155 288.270 168.470 ;
        RECT 282.385 168.135 282.765 168.155 ;
        RECT 287.885 168.135 288.265 168.155 ;
        RECT 291.885 168.135 292.265 168.515 ;
        RECT 295.885 168.135 296.265 168.515 ;
        RECT 301.595 168.435 303.335 168.725 ;
        RECT 305.385 168.385 306.585 168.675 ;
        RECT 308.095 168.345 310.725 168.800 ;
        RECT 312.305 168.450 312.685 168.830 ;
        RECT 217.150 167.730 230.975 168.030 ;
        RECT 232.650 167.565 248.660 167.940 ;
        RECT 266.475 167.510 287.250 167.885 ;
        RECT 217.155 166.985 235.575 167.285 ;
        RECT 237.020 166.975 264.330 167.315 ;
        RECT 216.635 166.270 223.895 166.570 ;
        RECT 5.325 165.650 9.450 165.920 ;
        RECT 36.285 165.845 54.955 165.855 ;
        RECT 36.285 165.800 66.305 165.845 ;
        RECT 36.285 165.790 93.545 165.800 ;
        RECT 36.285 165.535 102.550 165.790 ;
        RECT 201.690 165.650 205.815 165.920 ;
        RECT 217.190 165.735 221.275 166.005 ;
        RECT 227.595 165.970 231.345 166.245 ;
        RECT 232.650 166.210 258.880 166.600 ;
        RECT 265.505 166.155 297.470 166.545 ;
        RECT 310.280 165.915 313.410 166.190 ;
        RECT 314.155 166.155 314.535 173.315 ;
        RECT 363.900 171.185 365.100 171.565 ;
        RECT 315.395 170.855 322.135 171.155 ;
        RECT 366.855 170.970 369.130 171.480 ;
        RECT 371.755 170.970 374.055 171.480 ;
        RECT 376.350 170.970 378.630 171.480 ;
        RECT 383.425 171.285 384.660 171.665 ;
        RECT 315.985 169.060 319.440 169.500 ;
        RECT 322.445 168.900 322.825 169.280 ;
        RECT 363.900 168.885 367.160 169.265 ;
        RECT 367.900 168.885 371.160 169.265 ;
        RECT 377.400 168.885 380.660 169.265 ;
        RECT 381.400 168.885 384.660 169.265 ;
        RECT 320.845 168.385 322.045 168.675 ;
        RECT 327.765 168.450 328.145 168.830 ;
        RECT 314.800 167.675 330.720 167.975 ;
        RECT 315.335 166.930 332.280 167.230 ;
        RECT 364.565 166.970 390.860 167.310 ;
        RECT 396.950 166.160 397.330 173.320 ;
        RECT 398.780 169.105 402.155 169.505 ;
        RECT 402.525 168.865 402.905 169.245 ;
        RECT 405.240 168.905 405.620 169.285 ;
        RECT 409.425 168.855 409.805 169.235 ;
        RECT 399.850 168.440 401.590 168.730 ;
        RECT 403.640 168.390 404.840 168.680 ;
        RECT 406.350 168.360 408.960 168.785 ;
        RECT 410.560 168.455 410.940 168.835 ;
        RECT 398.095 167.680 411.660 167.995 ;
        RECT 398.090 166.935 411.650 167.235 ;
        RECT 398.110 166.220 404.835 166.520 ;
        RECT 408.535 165.920 411.640 166.195 ;
        RECT 412.410 166.160 412.790 173.320 ;
        RECT 468.860 173.265 525.215 173.320 ;
        RECT 429.050 172.280 466.600 172.335 ;
        RECT 429.050 172.050 494.620 172.280 ;
        RECT 465.845 171.995 494.620 172.050 ;
        RECT 496.290 171.975 502.995 172.275 ;
        RECT 430.560 171.140 432.015 171.520 ;
        RECT 432.755 171.140 433.955 171.520 ;
        RECT 435.710 170.925 437.985 171.435 ;
        RECT 440.610 170.925 442.910 171.435 ;
        RECT 445.205 170.925 447.485 171.435 ;
        RECT 452.280 171.240 453.515 171.620 ;
        RECT 454.255 171.240 455.535 171.620 ;
        RECT 469.150 171.085 470.605 171.465 ;
        RECT 453.695 170.885 454.075 170.920 ;
        RECT 432.195 170.780 432.575 170.820 ;
        RECT 432.125 170.475 434.960 170.780 ;
        RECT 450.940 170.575 454.075 170.885 ;
        RECT 474.300 170.870 476.575 171.380 ;
        RECT 479.200 170.870 481.500 171.380 ;
        RECT 483.795 170.870 486.075 171.380 ;
        RECT 492.845 171.185 494.125 171.565 ;
        RECT 492.285 170.830 492.665 170.865 ;
        RECT 470.785 170.725 471.165 170.765 ;
        RECT 453.695 170.540 454.075 170.575 ;
        RECT 432.195 170.440 432.575 170.475 ;
        RECT 470.715 170.420 473.550 170.725 ;
        RECT 489.530 170.520 492.665 170.830 ;
        RECT 492.285 170.485 492.665 170.520 ;
        RECT 470.785 170.385 471.165 170.420 ;
        RECT 414.240 169.065 417.645 169.505 ;
        RECT 417.985 168.865 418.365 169.245 ;
        RECT 420.700 168.905 421.080 169.285 ;
        RECT 424.885 168.855 425.265 169.235 ;
        RECT 430.720 168.840 432.015 169.220 ;
        RECT 432.755 168.840 436.015 169.220 ;
        RECT 436.755 168.840 440.015 169.220 ;
        RECT 440.755 168.840 441.940 169.220 ;
        RECT 444.205 168.840 445.515 169.220 ;
        RECT 446.255 168.840 449.515 169.220 ;
        RECT 450.255 168.840 453.515 169.220 ;
        RECT 454.255 168.840 455.270 169.220 ;
        RECT 415.310 168.440 417.050 168.730 ;
        RECT 419.100 168.390 420.300 168.680 ;
        RECT 421.810 168.360 424.405 168.735 ;
        RECT 426.020 168.455 426.400 168.835 ;
        RECT 469.310 168.785 470.605 169.165 ;
        RECT 475.345 168.785 478.605 169.165 ;
        RECT 479.345 168.785 480.530 169.165 ;
        RECT 482.795 168.785 484.105 169.165 ;
        RECT 484.845 168.785 488.105 169.165 ;
        RECT 492.845 168.785 493.860 169.165 ;
        RECT 496.925 169.030 500.340 169.450 ;
        RECT 500.670 168.810 501.050 169.190 ;
        RECT 503.385 168.850 503.765 169.230 ;
        RECT 507.570 168.800 507.950 169.180 ;
        RECT 432.195 168.140 432.575 168.520 ;
        RECT 436.195 168.140 436.575 168.520 ;
        RECT 440.195 168.475 440.575 168.520 ;
        RECT 445.695 168.475 446.075 168.520 ;
        RECT 440.145 168.160 446.080 168.475 ;
        RECT 440.195 168.140 440.575 168.160 ;
        RECT 445.695 168.140 446.075 168.160 ;
        RECT 449.695 168.140 450.075 168.520 ;
        RECT 453.695 168.140 454.075 168.520 ;
        RECT 470.785 168.085 471.165 168.465 ;
        RECT 474.785 168.085 475.165 168.465 ;
        RECT 478.785 168.420 479.165 168.465 ;
        RECT 484.285 168.420 484.665 168.465 ;
        RECT 478.735 168.105 484.670 168.420 ;
        RECT 478.785 168.085 479.165 168.105 ;
        RECT 484.285 168.085 484.665 168.105 ;
        RECT 488.285 168.085 488.665 168.465 ;
        RECT 492.285 168.085 492.665 168.465 ;
        RECT 497.995 168.385 499.735 168.675 ;
        RECT 501.785 168.335 502.985 168.625 ;
        RECT 504.495 168.295 507.125 168.750 ;
        RECT 508.705 168.400 509.085 168.780 ;
        RECT 413.550 167.680 427.375 167.980 ;
        RECT 429.050 167.515 445.060 167.890 ;
        RECT 462.875 167.460 483.650 167.835 ;
        RECT 413.555 166.935 431.975 167.235 ;
        RECT 433.420 166.925 460.730 167.265 ;
        RECT 413.035 166.220 420.295 166.520 ;
        RECT 232.650 165.845 251.320 165.855 ;
        RECT 232.650 165.800 262.670 165.845 ;
        RECT 232.650 165.790 289.910 165.800 ;
        RECT 232.650 165.535 298.915 165.790 ;
        RECT 398.090 165.600 402.215 165.870 ;
        RECT 413.590 165.685 417.675 165.955 ;
        RECT 423.995 165.920 427.745 166.195 ;
        RECT 429.050 166.160 455.280 166.550 ;
        RECT 461.905 166.105 493.870 166.495 ;
        RECT 506.680 165.865 509.810 166.140 ;
        RECT 510.555 166.105 510.935 173.265 ;
        RECT 560.220 171.230 561.420 171.610 ;
        RECT 511.795 170.805 518.535 171.105 ;
        RECT 563.175 171.015 565.450 171.525 ;
        RECT 568.075 171.015 570.375 171.525 ;
        RECT 572.670 171.015 574.950 171.525 ;
        RECT 579.745 171.330 580.980 171.710 ;
        RECT 512.385 169.010 515.840 169.450 ;
        RECT 518.845 168.850 519.225 169.230 ;
        RECT 560.220 168.930 563.480 169.310 ;
        RECT 564.220 168.930 567.480 169.310 ;
        RECT 573.720 168.930 576.980 169.310 ;
        RECT 577.720 168.930 580.980 169.310 ;
        RECT 517.245 168.335 518.445 168.625 ;
        RECT 524.165 168.400 524.545 168.780 ;
        RECT 511.200 167.625 527.120 167.925 ;
        RECT 511.735 166.880 528.680 167.180 ;
        RECT 560.885 167.015 587.180 167.355 ;
        RECT 593.325 166.195 593.705 173.355 ;
        RECT 595.155 169.140 598.530 169.540 ;
        RECT 598.900 168.900 599.280 169.280 ;
        RECT 601.615 168.940 601.995 169.320 ;
        RECT 605.800 168.890 606.180 169.270 ;
        RECT 596.225 168.475 597.965 168.765 ;
        RECT 600.015 168.425 601.215 168.715 ;
        RECT 602.725 168.395 605.335 168.820 ;
        RECT 606.935 168.490 607.315 168.870 ;
        RECT 594.470 167.715 608.035 168.030 ;
        RECT 594.465 166.970 608.025 167.270 ;
        RECT 594.485 166.255 601.210 166.555 ;
        RECT 604.910 165.955 608.015 166.230 ;
        RECT 608.785 166.195 609.165 173.355 ;
        RECT 665.235 173.300 721.590 173.355 ;
        RECT 625.425 172.315 662.975 172.370 ;
        RECT 625.425 172.085 690.995 172.315 ;
        RECT 662.220 172.030 690.995 172.085 ;
        RECT 692.665 172.010 699.370 172.310 ;
        RECT 626.935 171.175 628.390 171.555 ;
        RECT 629.130 171.175 630.330 171.555 ;
        RECT 632.085 170.960 634.360 171.470 ;
        RECT 636.985 170.960 639.285 171.470 ;
        RECT 641.580 170.960 643.860 171.470 ;
        RECT 648.655 171.275 649.890 171.655 ;
        RECT 650.630 171.275 651.910 171.655 ;
        RECT 665.525 171.120 666.980 171.500 ;
        RECT 650.070 170.920 650.450 170.955 ;
        RECT 628.570 170.815 628.950 170.855 ;
        RECT 628.500 170.510 631.335 170.815 ;
        RECT 647.315 170.610 650.450 170.920 ;
        RECT 670.675 170.905 672.950 171.415 ;
        RECT 675.575 170.905 677.875 171.415 ;
        RECT 680.170 170.905 682.450 171.415 ;
        RECT 689.220 171.220 690.500 171.600 ;
        RECT 688.660 170.865 689.040 170.900 ;
        RECT 667.160 170.760 667.540 170.800 ;
        RECT 650.070 170.575 650.450 170.610 ;
        RECT 628.570 170.475 628.950 170.510 ;
        RECT 667.090 170.455 669.925 170.760 ;
        RECT 685.905 170.555 689.040 170.865 ;
        RECT 688.660 170.520 689.040 170.555 ;
        RECT 667.160 170.420 667.540 170.455 ;
        RECT 610.615 169.100 614.020 169.540 ;
        RECT 614.360 168.900 614.740 169.280 ;
        RECT 617.075 168.940 617.455 169.320 ;
        RECT 621.260 168.890 621.640 169.270 ;
        RECT 627.095 168.875 628.390 169.255 ;
        RECT 629.130 168.875 632.390 169.255 ;
        RECT 633.130 168.875 636.390 169.255 ;
        RECT 637.130 168.875 638.315 169.255 ;
        RECT 640.580 168.875 641.890 169.255 ;
        RECT 642.630 168.875 645.890 169.255 ;
        RECT 646.630 168.875 649.890 169.255 ;
        RECT 650.630 168.875 651.645 169.255 ;
        RECT 611.685 168.475 613.425 168.765 ;
        RECT 615.475 168.425 616.675 168.715 ;
        RECT 618.185 168.395 620.780 168.770 ;
        RECT 622.395 168.490 622.775 168.870 ;
        RECT 665.685 168.820 666.980 169.200 ;
        RECT 671.720 168.820 674.980 169.200 ;
        RECT 675.720 168.820 676.905 169.200 ;
        RECT 679.170 168.820 680.480 169.200 ;
        RECT 681.220 168.820 684.480 169.200 ;
        RECT 689.220 168.820 690.235 169.200 ;
        RECT 693.300 169.065 696.715 169.485 ;
        RECT 697.045 168.845 697.425 169.225 ;
        RECT 699.760 168.885 700.140 169.265 ;
        RECT 703.945 168.835 704.325 169.215 ;
        RECT 628.570 168.175 628.950 168.555 ;
        RECT 632.570 168.175 632.950 168.555 ;
        RECT 636.570 168.510 636.950 168.555 ;
        RECT 642.070 168.510 642.450 168.555 ;
        RECT 636.520 168.195 642.455 168.510 ;
        RECT 636.570 168.175 636.950 168.195 ;
        RECT 642.070 168.175 642.450 168.195 ;
        RECT 646.070 168.175 646.450 168.555 ;
        RECT 650.070 168.175 650.450 168.555 ;
        RECT 667.160 168.120 667.540 168.500 ;
        RECT 671.160 168.120 671.540 168.500 ;
        RECT 675.160 168.455 675.540 168.500 ;
        RECT 680.660 168.455 681.040 168.500 ;
        RECT 675.110 168.140 681.045 168.455 ;
        RECT 675.160 168.120 675.540 168.140 ;
        RECT 680.660 168.120 681.040 168.140 ;
        RECT 684.660 168.120 685.040 168.500 ;
        RECT 688.660 168.120 689.040 168.500 ;
        RECT 694.370 168.420 696.110 168.710 ;
        RECT 698.160 168.370 699.360 168.660 ;
        RECT 700.870 168.330 703.500 168.785 ;
        RECT 705.080 168.435 705.460 168.815 ;
        RECT 609.925 167.715 623.750 168.015 ;
        RECT 625.425 167.550 641.435 167.925 ;
        RECT 659.250 167.495 680.025 167.870 ;
        RECT 609.930 166.970 628.350 167.270 ;
        RECT 629.795 166.960 657.105 167.300 ;
        RECT 609.410 166.255 616.670 166.555 ;
        RECT 429.050 165.795 447.720 165.805 ;
        RECT 429.050 165.750 459.070 165.795 ;
        RECT 429.050 165.740 486.310 165.750 ;
        RECT 65.985 165.480 102.550 165.535 ;
        RECT 262.350 165.480 298.915 165.535 ;
        RECT 429.050 165.485 495.315 165.740 ;
        RECT 594.465 165.635 598.590 165.905 ;
        RECT 609.965 165.720 614.050 165.990 ;
        RECT 620.370 165.955 624.120 166.230 ;
        RECT 625.425 166.195 651.655 166.585 ;
        RECT 658.280 166.140 690.245 166.530 ;
        RECT 703.055 165.900 706.185 166.175 ;
        RECT 706.930 166.140 707.310 173.300 ;
        RECT 756.585 171.235 757.785 171.615 ;
        RECT 708.170 170.840 714.910 171.140 ;
        RECT 759.540 171.020 761.815 171.530 ;
        RECT 764.440 171.020 766.740 171.530 ;
        RECT 769.035 171.020 771.315 171.530 ;
        RECT 776.110 171.335 777.345 171.715 ;
        RECT 708.760 169.045 712.215 169.485 ;
        RECT 715.220 168.885 715.600 169.265 ;
        RECT 756.585 168.935 759.845 169.315 ;
        RECT 760.585 168.935 763.845 169.315 ;
        RECT 770.085 168.935 773.345 169.315 ;
        RECT 774.085 168.935 777.345 169.315 ;
        RECT 713.620 168.370 714.820 168.660 ;
        RECT 720.540 168.435 720.920 168.815 ;
        RECT 707.575 167.660 723.495 167.960 ;
        RECT 708.110 166.915 725.055 167.215 ;
        RECT 757.250 167.020 783.545 167.360 ;
        RECT 789.665 166.195 790.045 173.355 ;
        RECT 791.495 169.140 794.870 169.540 ;
        RECT 795.240 168.900 795.620 169.280 ;
        RECT 797.955 168.940 798.335 169.320 ;
        RECT 802.140 168.890 802.520 169.270 ;
        RECT 792.565 168.475 794.305 168.765 ;
        RECT 796.355 168.425 797.555 168.715 ;
        RECT 799.065 168.395 801.675 168.820 ;
        RECT 803.275 168.490 803.655 168.870 ;
        RECT 790.810 167.715 804.375 168.030 ;
        RECT 790.805 166.970 804.365 167.270 ;
        RECT 790.825 166.255 797.550 166.555 ;
        RECT 801.250 165.955 804.355 166.230 ;
        RECT 805.125 166.195 805.505 173.355 ;
        RECT 861.575 173.300 917.930 173.355 ;
        RECT 821.765 172.315 859.315 172.370 ;
        RECT 821.765 172.085 887.335 172.315 ;
        RECT 858.560 172.030 887.335 172.085 ;
        RECT 889.005 172.010 895.710 172.310 ;
        RECT 823.275 171.175 824.730 171.555 ;
        RECT 825.470 171.175 826.670 171.555 ;
        RECT 828.425 170.960 830.700 171.470 ;
        RECT 833.325 170.960 835.625 171.470 ;
        RECT 837.920 170.960 840.200 171.470 ;
        RECT 844.995 171.275 846.230 171.655 ;
        RECT 846.970 171.275 848.250 171.655 ;
        RECT 861.865 171.120 863.320 171.500 ;
        RECT 846.410 170.920 846.790 170.955 ;
        RECT 824.910 170.815 825.290 170.855 ;
        RECT 824.840 170.510 827.675 170.815 ;
        RECT 843.655 170.610 846.790 170.920 ;
        RECT 867.015 170.905 869.290 171.415 ;
        RECT 871.915 170.905 874.215 171.415 ;
        RECT 876.510 170.905 878.790 171.415 ;
        RECT 885.560 171.220 886.840 171.600 ;
        RECT 885.000 170.865 885.380 170.900 ;
        RECT 863.500 170.760 863.880 170.800 ;
        RECT 846.410 170.575 846.790 170.610 ;
        RECT 824.910 170.475 825.290 170.510 ;
        RECT 863.430 170.455 866.265 170.760 ;
        RECT 882.245 170.555 885.380 170.865 ;
        RECT 885.000 170.520 885.380 170.555 ;
        RECT 863.500 170.420 863.880 170.455 ;
        RECT 806.955 169.100 810.360 169.540 ;
        RECT 810.700 168.900 811.080 169.280 ;
        RECT 813.415 168.940 813.795 169.320 ;
        RECT 817.600 168.890 817.980 169.270 ;
        RECT 823.435 168.875 824.730 169.255 ;
        RECT 825.470 168.875 828.730 169.255 ;
        RECT 829.470 168.875 832.730 169.255 ;
        RECT 833.470 168.875 834.655 169.255 ;
        RECT 836.920 168.875 838.230 169.255 ;
        RECT 838.970 168.875 842.230 169.255 ;
        RECT 842.970 168.875 846.230 169.255 ;
        RECT 846.970 168.875 847.985 169.255 ;
        RECT 808.025 168.475 809.765 168.765 ;
        RECT 811.815 168.425 813.015 168.715 ;
        RECT 814.525 168.395 817.120 168.770 ;
        RECT 818.735 168.490 819.115 168.870 ;
        RECT 862.025 168.820 863.320 169.200 ;
        RECT 868.060 168.820 871.320 169.200 ;
        RECT 872.060 168.820 873.245 169.200 ;
        RECT 875.510 168.820 876.820 169.200 ;
        RECT 877.560 168.820 880.820 169.200 ;
        RECT 885.560 168.820 886.575 169.200 ;
        RECT 889.640 169.065 893.055 169.485 ;
        RECT 893.385 168.845 893.765 169.225 ;
        RECT 896.100 168.885 896.480 169.265 ;
        RECT 900.285 168.835 900.665 169.215 ;
        RECT 824.910 168.175 825.290 168.555 ;
        RECT 828.910 168.175 829.290 168.555 ;
        RECT 832.910 168.510 833.290 168.555 ;
        RECT 838.410 168.510 838.790 168.555 ;
        RECT 832.860 168.195 838.795 168.510 ;
        RECT 832.910 168.175 833.290 168.195 ;
        RECT 838.410 168.175 838.790 168.195 ;
        RECT 842.410 168.175 842.790 168.555 ;
        RECT 846.410 168.175 846.790 168.555 ;
        RECT 863.500 168.120 863.880 168.500 ;
        RECT 867.500 168.120 867.880 168.500 ;
        RECT 871.500 168.455 871.880 168.500 ;
        RECT 877.000 168.455 877.380 168.500 ;
        RECT 871.450 168.140 877.385 168.455 ;
        RECT 871.500 168.120 871.880 168.140 ;
        RECT 877.000 168.120 877.380 168.140 ;
        RECT 881.000 168.120 881.380 168.500 ;
        RECT 885.000 168.120 885.380 168.500 ;
        RECT 890.710 168.420 892.450 168.710 ;
        RECT 894.500 168.370 895.700 168.660 ;
        RECT 897.210 168.330 899.840 168.785 ;
        RECT 901.420 168.435 901.800 168.815 ;
        RECT 806.265 167.715 820.090 168.015 ;
        RECT 821.765 167.550 837.775 167.925 ;
        RECT 855.590 167.495 876.365 167.870 ;
        RECT 806.270 166.970 824.690 167.270 ;
        RECT 826.135 166.960 853.445 167.300 ;
        RECT 805.750 166.255 813.010 166.555 ;
        RECT 625.425 165.830 644.095 165.840 ;
        RECT 625.425 165.785 655.445 165.830 ;
        RECT 625.425 165.775 682.685 165.785 ;
        RECT 625.425 165.520 691.690 165.775 ;
        RECT 790.805 165.635 794.930 165.905 ;
        RECT 806.305 165.720 810.390 165.990 ;
        RECT 816.710 165.955 820.460 166.230 ;
        RECT 821.765 166.195 847.995 166.585 ;
        RECT 854.620 166.140 886.585 166.530 ;
        RECT 899.395 165.900 902.525 166.175 ;
        RECT 903.270 166.140 903.650 173.300 ;
        RECT 952.970 171.220 954.170 171.600 ;
        RECT 904.510 170.840 911.250 171.140 ;
        RECT 955.925 171.005 958.200 171.515 ;
        RECT 960.825 171.005 963.125 171.515 ;
        RECT 965.420 171.005 967.700 171.515 ;
        RECT 972.495 171.320 973.730 171.700 ;
        RECT 905.100 169.045 908.555 169.485 ;
        RECT 911.560 168.885 911.940 169.265 ;
        RECT 952.970 168.920 956.230 169.300 ;
        RECT 956.970 168.920 960.230 169.300 ;
        RECT 966.470 168.920 969.730 169.300 ;
        RECT 970.470 168.920 973.730 169.300 ;
        RECT 909.960 168.370 911.160 168.660 ;
        RECT 916.880 168.435 917.260 168.815 ;
        RECT 903.915 167.660 919.835 167.960 ;
        RECT 904.450 166.915 921.395 167.215 ;
        RECT 953.635 167.005 979.930 167.345 ;
        RECT 986.005 166.195 986.385 173.355 ;
        RECT 987.835 169.140 991.210 169.540 ;
        RECT 991.580 168.900 991.960 169.280 ;
        RECT 994.295 168.940 994.675 169.320 ;
        RECT 998.480 168.890 998.860 169.270 ;
        RECT 988.905 168.475 990.645 168.765 ;
        RECT 992.695 168.425 993.895 168.715 ;
        RECT 995.405 168.395 998.015 168.820 ;
        RECT 999.615 168.490 999.995 168.870 ;
        RECT 987.150 167.715 1000.715 168.030 ;
        RECT 987.145 166.970 1000.705 167.270 ;
        RECT 987.165 166.255 993.890 166.555 ;
        RECT 997.590 165.955 1000.695 166.230 ;
        RECT 1001.465 166.195 1001.845 173.355 ;
        RECT 1057.915 173.300 1114.270 173.355 ;
        RECT 1018.105 172.315 1055.655 172.370 ;
        RECT 1018.105 172.085 1083.675 172.315 ;
        RECT 1054.900 172.030 1083.675 172.085 ;
        RECT 1085.345 172.010 1092.050 172.310 ;
        RECT 1019.615 171.175 1021.070 171.555 ;
        RECT 1021.810 171.175 1023.010 171.555 ;
        RECT 1024.765 170.960 1027.040 171.470 ;
        RECT 1029.665 170.960 1031.965 171.470 ;
        RECT 1034.260 170.960 1036.540 171.470 ;
        RECT 1041.335 171.275 1042.570 171.655 ;
        RECT 1043.310 171.275 1044.590 171.655 ;
        RECT 1058.205 171.120 1059.660 171.500 ;
        RECT 1042.750 170.920 1043.130 170.955 ;
        RECT 1021.250 170.815 1021.630 170.855 ;
        RECT 1021.180 170.510 1024.015 170.815 ;
        RECT 1039.995 170.610 1043.130 170.920 ;
        RECT 1063.355 170.905 1065.630 171.415 ;
        RECT 1068.255 170.905 1070.555 171.415 ;
        RECT 1072.850 170.905 1075.130 171.415 ;
        RECT 1081.900 171.220 1083.180 171.600 ;
        RECT 1081.340 170.865 1081.720 170.900 ;
        RECT 1059.840 170.760 1060.220 170.800 ;
        RECT 1042.750 170.575 1043.130 170.610 ;
        RECT 1021.250 170.475 1021.630 170.510 ;
        RECT 1059.770 170.455 1062.605 170.760 ;
        RECT 1078.585 170.555 1081.720 170.865 ;
        RECT 1081.340 170.520 1081.720 170.555 ;
        RECT 1059.840 170.420 1060.220 170.455 ;
        RECT 1003.295 169.100 1006.700 169.540 ;
        RECT 1007.040 168.900 1007.420 169.280 ;
        RECT 1009.755 168.940 1010.135 169.320 ;
        RECT 1013.940 168.890 1014.320 169.270 ;
        RECT 1019.775 168.875 1021.070 169.255 ;
        RECT 1021.810 168.875 1025.070 169.255 ;
        RECT 1025.810 168.875 1029.070 169.255 ;
        RECT 1029.810 168.875 1030.995 169.255 ;
        RECT 1033.260 168.875 1034.570 169.255 ;
        RECT 1035.310 168.875 1038.570 169.255 ;
        RECT 1039.310 168.875 1042.570 169.255 ;
        RECT 1043.310 168.875 1044.325 169.255 ;
        RECT 1004.365 168.475 1006.105 168.765 ;
        RECT 1008.155 168.425 1009.355 168.715 ;
        RECT 1010.865 168.395 1013.460 168.770 ;
        RECT 1015.075 168.490 1015.455 168.870 ;
        RECT 1058.365 168.820 1059.660 169.200 ;
        RECT 1064.400 168.820 1067.660 169.200 ;
        RECT 1068.400 168.820 1069.585 169.200 ;
        RECT 1071.850 168.820 1073.160 169.200 ;
        RECT 1073.900 168.820 1077.160 169.200 ;
        RECT 1081.900 168.820 1082.915 169.200 ;
        RECT 1085.980 169.065 1089.395 169.485 ;
        RECT 1089.725 168.845 1090.105 169.225 ;
        RECT 1092.440 168.885 1092.820 169.265 ;
        RECT 1096.625 168.835 1097.005 169.215 ;
        RECT 1021.250 168.175 1021.630 168.555 ;
        RECT 1025.250 168.175 1025.630 168.555 ;
        RECT 1029.250 168.510 1029.630 168.555 ;
        RECT 1034.750 168.510 1035.130 168.555 ;
        RECT 1029.200 168.195 1035.135 168.510 ;
        RECT 1029.250 168.175 1029.630 168.195 ;
        RECT 1034.750 168.175 1035.130 168.195 ;
        RECT 1038.750 168.175 1039.130 168.555 ;
        RECT 1042.750 168.175 1043.130 168.555 ;
        RECT 1059.840 168.120 1060.220 168.500 ;
        RECT 1063.840 168.120 1064.220 168.500 ;
        RECT 1067.840 168.455 1068.220 168.500 ;
        RECT 1073.340 168.455 1073.720 168.500 ;
        RECT 1067.790 168.140 1073.725 168.455 ;
        RECT 1067.840 168.120 1068.220 168.140 ;
        RECT 1073.340 168.120 1073.720 168.140 ;
        RECT 1077.340 168.120 1077.720 168.500 ;
        RECT 1081.340 168.120 1081.720 168.500 ;
        RECT 1087.050 168.420 1088.790 168.710 ;
        RECT 1090.840 168.370 1092.040 168.660 ;
        RECT 1093.550 168.330 1096.180 168.785 ;
        RECT 1097.760 168.435 1098.140 168.815 ;
        RECT 1002.605 167.715 1016.430 168.015 ;
        RECT 1018.105 167.550 1034.115 167.925 ;
        RECT 1051.930 167.495 1072.705 167.870 ;
        RECT 1002.610 166.970 1021.030 167.270 ;
        RECT 1022.475 166.960 1049.785 167.300 ;
        RECT 1002.090 166.255 1009.350 166.555 ;
        RECT 821.765 165.830 840.435 165.840 ;
        RECT 821.765 165.785 851.785 165.830 ;
        RECT 821.765 165.775 879.025 165.785 ;
        RECT 821.765 165.520 888.030 165.775 ;
        RECT 987.145 165.635 991.270 165.905 ;
        RECT 1002.645 165.720 1006.730 165.990 ;
        RECT 1013.050 165.955 1016.800 166.230 ;
        RECT 1018.105 166.195 1044.335 166.585 ;
        RECT 1050.960 166.140 1082.925 166.530 ;
        RECT 1095.735 165.900 1098.865 166.175 ;
        RECT 1099.610 166.140 1099.990 173.300 ;
        RECT 1149.295 171.225 1150.495 171.605 ;
        RECT 1100.850 170.840 1107.590 171.140 ;
        RECT 1152.250 171.010 1154.525 171.520 ;
        RECT 1157.150 171.010 1159.450 171.520 ;
        RECT 1161.745 171.010 1164.025 171.520 ;
        RECT 1168.820 171.325 1170.055 171.705 ;
        RECT 1101.440 169.045 1104.895 169.485 ;
        RECT 1107.900 168.885 1108.280 169.265 ;
        RECT 1149.295 168.925 1152.555 169.305 ;
        RECT 1153.295 168.925 1156.555 169.305 ;
        RECT 1162.795 168.925 1166.055 169.305 ;
        RECT 1166.795 168.925 1170.055 169.305 ;
        RECT 1106.300 168.370 1107.500 168.660 ;
        RECT 1113.220 168.435 1113.600 168.815 ;
        RECT 1100.255 167.660 1116.175 167.960 ;
        RECT 1100.790 166.915 1117.735 167.215 ;
        RECT 1149.960 167.010 1176.255 167.350 ;
        RECT 1182.345 166.195 1182.725 173.355 ;
        RECT 1184.175 169.140 1187.550 169.540 ;
        RECT 1187.920 168.900 1188.300 169.280 ;
        RECT 1190.635 168.940 1191.015 169.320 ;
        RECT 1194.820 168.890 1195.200 169.270 ;
        RECT 1185.245 168.475 1186.985 168.765 ;
        RECT 1189.035 168.425 1190.235 168.715 ;
        RECT 1191.745 168.395 1194.355 168.820 ;
        RECT 1195.955 168.490 1196.335 168.870 ;
        RECT 1183.490 167.715 1197.055 168.030 ;
        RECT 1183.485 166.970 1197.045 167.270 ;
        RECT 1183.505 166.255 1190.230 166.555 ;
        RECT 1193.930 165.955 1197.035 166.230 ;
        RECT 1197.805 166.195 1198.185 173.355 ;
        RECT 1254.255 173.300 1310.610 173.355 ;
        RECT 1214.445 172.315 1251.995 172.370 ;
        RECT 1214.445 172.085 1280.015 172.315 ;
        RECT 1251.240 172.030 1280.015 172.085 ;
        RECT 1281.685 172.010 1288.390 172.310 ;
        RECT 1215.955 171.175 1217.410 171.555 ;
        RECT 1218.150 171.175 1219.350 171.555 ;
        RECT 1221.105 170.960 1223.380 171.470 ;
        RECT 1226.005 170.960 1228.305 171.470 ;
        RECT 1230.600 170.960 1232.880 171.470 ;
        RECT 1237.675 171.275 1238.910 171.655 ;
        RECT 1239.650 171.275 1240.930 171.655 ;
        RECT 1254.545 171.120 1256.000 171.500 ;
        RECT 1256.740 171.120 1257.940 171.500 ;
        RECT 1239.090 170.920 1239.470 170.955 ;
        RECT 1217.590 170.815 1217.970 170.855 ;
        RECT 1217.520 170.510 1220.355 170.815 ;
        RECT 1236.335 170.610 1239.470 170.920 ;
        RECT 1259.695 170.905 1261.970 171.415 ;
        RECT 1264.595 170.905 1266.895 171.415 ;
        RECT 1269.190 170.905 1271.470 171.415 ;
        RECT 1276.265 171.220 1277.500 171.600 ;
        RECT 1278.240 171.220 1279.520 171.600 ;
        RECT 1277.680 170.865 1278.060 170.900 ;
        RECT 1256.180 170.760 1256.560 170.800 ;
        RECT 1239.090 170.575 1239.470 170.610 ;
        RECT 1217.590 170.475 1217.970 170.510 ;
        RECT 1256.110 170.455 1258.945 170.760 ;
        RECT 1274.925 170.555 1278.060 170.865 ;
        RECT 1277.680 170.520 1278.060 170.555 ;
        RECT 1256.180 170.420 1256.560 170.455 ;
        RECT 1199.635 169.100 1203.040 169.540 ;
        RECT 1203.380 168.900 1203.760 169.280 ;
        RECT 1206.095 168.940 1206.475 169.320 ;
        RECT 1210.280 168.890 1210.660 169.270 ;
        RECT 1216.115 168.875 1217.410 169.255 ;
        RECT 1218.150 168.875 1221.410 169.255 ;
        RECT 1222.150 168.875 1225.410 169.255 ;
        RECT 1226.150 168.875 1227.335 169.255 ;
        RECT 1229.600 168.875 1230.910 169.255 ;
        RECT 1231.650 168.875 1234.910 169.255 ;
        RECT 1235.650 168.875 1238.910 169.255 ;
        RECT 1239.650 168.875 1240.665 169.255 ;
        RECT 1200.705 168.475 1202.445 168.765 ;
        RECT 1204.495 168.425 1205.695 168.715 ;
        RECT 1207.205 168.395 1209.800 168.770 ;
        RECT 1211.415 168.490 1211.795 168.870 ;
        RECT 1254.705 168.820 1256.000 169.200 ;
        RECT 1256.740 168.820 1260.000 169.200 ;
        RECT 1260.740 168.820 1264.000 169.200 ;
        RECT 1264.740 168.820 1265.925 169.200 ;
        RECT 1268.190 168.820 1269.500 169.200 ;
        RECT 1270.240 168.820 1273.500 169.200 ;
        RECT 1274.240 168.820 1277.500 169.200 ;
        RECT 1278.240 168.820 1279.255 169.200 ;
        RECT 1282.320 169.065 1285.735 169.485 ;
        RECT 1286.065 168.845 1286.445 169.225 ;
        RECT 1288.780 168.885 1289.160 169.265 ;
        RECT 1292.965 168.835 1293.345 169.215 ;
        RECT 1217.590 168.175 1217.970 168.555 ;
        RECT 1221.590 168.175 1221.970 168.555 ;
        RECT 1225.590 168.510 1225.970 168.555 ;
        RECT 1231.090 168.510 1231.470 168.555 ;
        RECT 1225.540 168.195 1231.475 168.510 ;
        RECT 1225.590 168.175 1225.970 168.195 ;
        RECT 1231.090 168.175 1231.470 168.195 ;
        RECT 1235.090 168.175 1235.470 168.555 ;
        RECT 1239.090 168.175 1239.470 168.555 ;
        RECT 1256.180 168.120 1256.560 168.500 ;
        RECT 1260.180 168.120 1260.560 168.500 ;
        RECT 1264.180 168.455 1264.560 168.500 ;
        RECT 1269.680 168.455 1270.060 168.500 ;
        RECT 1264.130 168.140 1270.065 168.455 ;
        RECT 1264.180 168.120 1264.560 168.140 ;
        RECT 1269.680 168.120 1270.060 168.140 ;
        RECT 1273.680 168.120 1274.060 168.500 ;
        RECT 1277.680 168.120 1278.060 168.500 ;
        RECT 1283.390 168.420 1285.130 168.710 ;
        RECT 1287.180 168.370 1288.380 168.660 ;
        RECT 1289.890 168.330 1292.520 168.785 ;
        RECT 1294.100 168.435 1294.480 168.815 ;
        RECT 1198.945 167.715 1212.770 168.015 ;
        RECT 1214.445 167.550 1230.455 167.925 ;
        RECT 1248.270 167.495 1269.045 167.870 ;
        RECT 1281.670 167.660 1295.285 167.960 ;
        RECT 1198.950 166.970 1217.370 167.270 ;
        RECT 1218.815 166.960 1246.125 167.300 ;
        RECT 1257.405 166.905 1279.960 167.245 ;
        RECT 1281.070 166.915 1295.715 167.215 ;
        RECT 1198.430 166.255 1205.690 166.555 ;
        RECT 1018.105 165.830 1036.775 165.840 ;
        RECT 1018.105 165.785 1048.125 165.830 ;
        RECT 1018.105 165.775 1075.365 165.785 ;
        RECT 1018.105 165.520 1084.370 165.775 ;
        RECT 1183.485 165.635 1187.610 165.905 ;
        RECT 1198.985 165.720 1203.070 165.990 ;
        RECT 1209.390 165.955 1213.140 166.230 ;
        RECT 1214.445 166.195 1240.675 166.585 ;
        RECT 1247.300 166.140 1279.265 166.530 ;
        RECT 1292.075 165.900 1295.205 166.175 ;
        RECT 1295.950 166.140 1296.330 173.300 ;
        RECT 1297.190 170.840 1303.930 171.140 ;
        RECT 1297.780 169.045 1301.235 169.485 ;
        RECT 1304.240 168.885 1304.620 169.265 ;
        RECT 1302.640 168.370 1303.840 168.660 ;
        RECT 1309.560 168.435 1309.940 168.815 ;
        RECT 1296.595 167.660 1312.515 167.960 ;
        RECT 1297.130 166.915 1314.075 167.215 ;
        RECT 1214.445 165.830 1233.115 165.840 ;
        RECT 1214.445 165.785 1244.465 165.830 ;
        RECT 1214.445 165.775 1271.705 165.785 ;
        RECT 1214.445 165.520 1280.710 165.775 ;
        RECT 458.750 165.430 495.315 165.485 ;
        RECT 655.125 165.465 691.690 165.520 ;
        RECT 851.465 165.465 888.030 165.520 ;
        RECT 1047.805 165.465 1084.370 165.520 ;
        RECT 1244.145 165.465 1280.710 165.520 ;
        RECT 6.560 165.075 10.690 165.375 ;
        RECT -59.600 164.300 -56.035 164.310 ;
        RECT -59.600 163.975 -55.240 164.300 ;
        RECT -9.275 164.055 -3.360 164.390 ;
        RECT -6.005 164.035 -3.360 164.055 ;
        RECT -56.195 163.965 -55.240 163.975 ;
        RECT -79.005 163.335 -75.705 163.715 ;
        RECT -75.005 163.335 -71.705 163.715 ;
        RECT -65.505 163.335 -62.205 163.715 ;
        RECT -61.505 163.335 -58.205 163.715 ;
        RECT -28.680 163.415 -25.380 163.795 ;
        RECT -24.680 163.415 -21.380 163.795 ;
        RECT -15.180 163.415 -11.880 163.795 ;
        RECT -11.180 163.415 -7.880 163.795 ;
        RECT -79.005 161.335 -77.720 161.715 ;
        RECT -59.690 161.335 -58.205 161.715 ;
        RECT -28.680 161.415 -27.395 161.795 ;
        RECT -9.365 161.415 -7.880 161.795 ;
        RECT -77.500 160.655 -75.980 161.015 ;
        RECT -27.175 160.735 -25.655 161.095 ;
        RECT -82.690 158.290 -56.035 159.190 ;
        RECT -32.365 158.370 -5.710 159.270 ;
        RECT 4.185 159.245 4.565 165.075 ;
        RECT 13.065 165.025 17.565 165.335 ;
        RECT 22.020 165.075 26.150 165.375 ;
        RECT 9.025 164.475 15.415 164.765 ;
        RECT 8.440 163.895 19.095 164.230 ;
        RECT 7.790 163.310 10.710 163.610 ;
        RECT 14.255 163.295 17.625 163.595 ;
        RECT 6.005 162.560 6.385 162.940 ;
        RECT 8.410 162.575 10.190 162.865 ;
        RECT 11.665 162.665 12.855 162.950 ;
        RECT 15.785 162.545 17.095 162.865 ;
        RECT 7.140 161.960 7.520 162.340 ;
        RECT 10.885 162.000 11.265 162.380 ;
        RECT 13.595 161.990 13.975 162.370 ;
        RECT 15.005 161.835 18.185 162.155 ;
        RECT 4.935 159.245 9.030 159.250 ;
        RECT 19.645 159.245 20.025 165.075 ;
        RECT 28.525 165.025 33.025 165.335 ;
        RECT 202.925 165.075 207.055 165.375 ;
        RECT 35.755 164.810 71.665 164.865 ;
        RECT 35.755 164.595 102.950 164.810 ;
        RECT 71.205 164.540 102.950 164.595 ;
        RECT 107.170 164.420 113.560 164.710 ;
        RECT 23.900 163.895 34.405 164.230 ;
        RECT 59.375 164.030 69.925 164.365 ;
        RECT 23.250 163.310 26.170 163.610 ;
        RECT 29.715 163.295 33.085 163.595 ;
        RECT 37.965 163.390 39.270 163.770 ;
        RECT 39.970 163.390 43.270 163.770 ;
        RECT 43.970 163.390 47.270 163.770 ;
        RECT 47.970 163.390 49.330 163.770 ;
        RECT 51.305 163.390 52.770 163.770 ;
        RECT 53.470 163.390 56.770 163.770 ;
        RECT 57.470 163.390 60.770 163.770 ;
        RECT 61.470 163.390 62.650 163.770 ;
        RECT 76.555 163.335 77.860 163.715 ;
        RECT 82.560 163.335 85.860 163.715 ;
        RECT 86.560 163.335 87.920 163.715 ;
        RECT 89.895 163.335 91.360 163.715 ;
        RECT 92.060 163.335 95.360 163.715 ;
        RECT 100.060 163.335 101.240 163.715 ;
        RECT 39.430 163.045 39.810 163.080 ;
        RECT 23.870 162.575 25.650 162.865 ;
        RECT 31.245 162.545 32.555 162.865 ;
        RECT 39.165 162.735 42.175 163.045 ;
        RECT 39.430 162.700 39.810 162.735 ;
        RECT 43.430 162.700 44.520 163.080 ;
        RECT 47.430 163.075 47.810 163.080 ;
        RECT 44.950 162.710 47.815 163.075 ;
        RECT 52.930 163.055 53.310 163.080 ;
        RECT 52.915 162.735 55.060 163.055 ;
        RECT 47.430 162.700 47.810 162.710 ;
        RECT 52.930 162.700 53.310 162.735 ;
        RECT 55.975 162.700 57.310 163.080 ;
        RECT 60.930 163.060 61.310 163.080 ;
        RECT 58.465 162.740 61.375 163.060 ;
        RECT 78.020 162.990 78.400 163.025 ;
        RECT 60.930 162.700 61.310 162.740 ;
        RECT 77.755 162.680 80.765 162.990 ;
        RECT 78.020 162.645 78.400 162.680 ;
        RECT 82.020 162.645 83.110 163.025 ;
        RECT 86.020 163.020 86.400 163.025 ;
        RECT 83.540 162.655 86.405 163.020 ;
        RECT 91.520 163.000 91.900 163.025 ;
        RECT 91.505 162.680 93.650 163.000 ;
        RECT 86.020 162.645 86.400 162.655 ;
        RECT 91.520 162.645 91.900 162.680 ;
        RECT 94.565 162.645 95.900 163.025 ;
        RECT 99.520 163.005 99.900 163.025 ;
        RECT 97.055 162.685 99.965 163.005 ;
        RECT 99.520 162.645 99.900 162.685 ;
        RECT 104.150 162.505 104.530 162.885 ;
        RECT 109.810 162.610 111.000 162.895 ;
        RECT 22.600 161.960 22.980 162.340 ;
        RECT 29.055 161.990 29.435 162.370 ;
        RECT 109.030 161.945 109.410 162.325 ;
        RECT 113.150 161.780 116.330 162.100 ;
        RECT 37.780 161.390 39.270 161.770 ;
        RECT 39.970 161.390 41.255 161.770 ;
        RECT 59.285 161.390 60.770 161.770 ;
        RECT 61.470 161.390 62.545 161.770 ;
        RECT 76.370 161.335 77.860 161.715 ;
        RECT 100.060 161.335 101.135 161.715 ;
        RECT 39.430 160.700 40.520 161.080 ;
        RECT 41.475 160.710 42.995 161.070 ;
        RECT 43.915 160.705 56.765 161.040 ;
        RECT 60.930 161.035 61.310 161.080 ;
        RECT 60.195 160.735 61.505 161.035 ;
        RECT 60.930 160.700 61.310 160.735 ;
        RECT 78.020 160.645 79.110 161.025 ;
        RECT 80.065 160.655 81.585 161.015 ;
        RECT 82.505 160.650 95.355 160.985 ;
        RECT 99.520 160.980 99.900 161.025 ;
        RECT 98.785 160.680 100.095 160.980 ;
        RECT 99.520 160.645 99.900 160.680 ;
        RECT 36.285 160.150 69.365 160.190 ;
        RECT 36.285 159.840 101.530 160.150 ;
        RECT 68.580 159.785 101.530 159.840 ;
        RECT 103.325 159.775 107.585 160.130 ;
        RECT 20.395 159.245 24.490 159.250 ;
        RECT 3.815 159.240 9.030 159.245 ;
        RECT 19.275 159.240 24.490 159.245 ;
        RECT 34.735 159.240 74.985 159.245 ;
        RECT 3.815 159.190 74.985 159.240 ;
        RECT 101.530 159.190 107.175 159.195 ;
        RECT 117.790 159.190 118.170 165.020 ;
        RECT 122.630 164.420 129.020 164.710 ;
        RECT 186.895 164.065 192.810 164.400 ;
        RECT 190.165 164.045 192.810 164.065 ;
        RECT 167.490 163.425 170.790 163.805 ;
        RECT 171.490 163.425 174.790 163.805 ;
        RECT 180.990 163.425 184.290 163.805 ;
        RECT 184.990 163.425 188.290 163.805 ;
        RECT 119.610 162.505 119.990 162.885 ;
        RECT 125.270 162.610 126.460 162.895 ;
        RECT 124.490 161.945 124.870 162.325 ;
        RECT 128.610 161.780 131.790 162.100 ;
        RECT 167.490 161.425 168.775 161.805 ;
        RECT 186.805 161.425 188.290 161.805 ;
        RECT 118.890 160.695 123.040 160.965 ;
        RECT 168.995 160.745 170.515 161.105 ;
        RECT 118.540 159.190 122.635 159.195 ;
        RECT 3.815 159.185 107.175 159.190 ;
        RECT 117.420 159.185 122.635 159.190 ;
        RECT 3.815 158.345 132.450 159.185 ;
        RECT 163.805 158.380 190.460 159.280 ;
        RECT 200.550 159.245 200.930 165.075 ;
        RECT 209.430 165.025 213.930 165.335 ;
        RECT 218.385 165.075 222.515 165.375 ;
        RECT 205.390 164.475 211.780 164.765 ;
        RECT 204.805 163.895 215.460 164.230 ;
        RECT 204.155 163.310 207.075 163.610 ;
        RECT 210.620 163.295 213.990 163.595 ;
        RECT 202.370 162.560 202.750 162.940 ;
        RECT 204.775 162.575 206.555 162.865 ;
        RECT 208.030 162.665 209.220 162.950 ;
        RECT 212.150 162.545 213.460 162.865 ;
        RECT 203.505 161.960 203.885 162.340 ;
        RECT 207.250 162.000 207.630 162.380 ;
        RECT 209.960 161.990 210.340 162.370 ;
        RECT 211.370 161.835 214.550 162.155 ;
        RECT 201.300 159.245 205.395 159.250 ;
        RECT 216.010 159.245 216.390 165.075 ;
        RECT 224.890 165.025 229.390 165.335 ;
        RECT 316.530 165.020 320.660 165.320 ;
        RECT 232.120 164.810 268.030 164.865 ;
        RECT 220.850 164.475 227.240 164.765 ;
        RECT 232.120 164.595 299.315 164.810 ;
        RECT 267.570 164.540 299.315 164.595 ;
        RECT 303.535 164.420 309.925 164.710 ;
        RECT 220.265 163.895 230.770 164.230 ;
        RECT 255.740 164.030 266.290 164.365 ;
        RECT 302.950 163.840 313.430 164.175 ;
        RECT 219.615 163.310 222.535 163.610 ;
        RECT 226.080 163.295 229.450 163.595 ;
        RECT 234.330 163.390 235.635 163.770 ;
        RECT 236.335 163.390 239.635 163.770 ;
        RECT 240.335 163.390 243.635 163.770 ;
        RECT 244.335 163.390 245.695 163.770 ;
        RECT 247.670 163.390 249.135 163.770 ;
        RECT 249.835 163.390 253.135 163.770 ;
        RECT 253.835 163.390 257.135 163.770 ;
        RECT 257.835 163.390 259.015 163.770 ;
        RECT 272.920 163.335 274.225 163.715 ;
        RECT 278.925 163.335 282.225 163.715 ;
        RECT 282.925 163.335 284.285 163.715 ;
        RECT 286.260 163.335 287.725 163.715 ;
        RECT 288.425 163.335 291.725 163.715 ;
        RECT 296.425 163.335 297.605 163.715 ;
        RECT 235.795 163.045 236.175 163.080 ;
        RECT 217.830 162.560 218.210 162.940 ;
        RECT 220.235 162.575 222.015 162.865 ;
        RECT 223.490 162.665 224.680 162.950 ;
        RECT 227.610 162.545 228.920 162.865 ;
        RECT 235.530 162.735 238.540 163.045 ;
        RECT 235.795 162.700 236.175 162.735 ;
        RECT 239.795 162.700 240.885 163.080 ;
        RECT 243.795 163.075 244.175 163.080 ;
        RECT 241.315 162.710 244.180 163.075 ;
        RECT 249.295 163.055 249.675 163.080 ;
        RECT 249.280 162.735 251.425 163.055 ;
        RECT 243.795 162.700 244.175 162.710 ;
        RECT 249.295 162.700 249.675 162.735 ;
        RECT 252.340 162.700 253.675 163.080 ;
        RECT 257.295 163.060 257.675 163.080 ;
        RECT 254.830 162.740 257.740 163.060 ;
        RECT 274.385 162.990 274.765 163.025 ;
        RECT 257.295 162.700 257.675 162.740 ;
        RECT 274.120 162.680 277.130 162.990 ;
        RECT 274.385 162.645 274.765 162.680 ;
        RECT 278.385 162.645 279.475 163.025 ;
        RECT 282.385 163.020 282.765 163.025 ;
        RECT 279.905 162.655 282.770 163.020 ;
        RECT 287.885 163.000 288.265 163.025 ;
        RECT 287.870 162.680 290.015 163.000 ;
        RECT 282.385 162.645 282.765 162.655 ;
        RECT 287.885 162.645 288.265 162.680 ;
        RECT 290.930 162.645 292.265 163.025 ;
        RECT 295.885 163.005 296.265 163.025 ;
        RECT 293.420 162.685 296.330 163.005 ;
        RECT 295.885 162.645 296.265 162.685 ;
        RECT 300.515 162.505 300.895 162.885 ;
        RECT 302.920 162.520 304.700 162.810 ;
        RECT 306.175 162.610 307.365 162.895 ;
        RECT 310.295 162.490 311.605 162.810 ;
        RECT 218.965 161.960 219.345 162.340 ;
        RECT 222.710 162.000 223.090 162.380 ;
        RECT 225.420 161.990 225.800 162.370 ;
        RECT 226.830 161.835 230.010 162.155 ;
        RECT 301.650 161.905 302.030 162.285 ;
        RECT 305.395 161.945 305.775 162.325 ;
        RECT 308.105 161.935 308.485 162.315 ;
        RECT 309.515 161.780 312.695 162.100 ;
        RECT 234.145 161.390 235.635 161.770 ;
        RECT 236.335 161.390 237.620 161.770 ;
        RECT 255.650 161.390 257.135 161.770 ;
        RECT 257.835 161.390 258.910 161.770 ;
        RECT 272.735 161.335 274.225 161.715 ;
        RECT 296.425 161.335 297.500 161.715 ;
        RECT 235.795 160.700 236.885 161.080 ;
        RECT 237.840 160.710 239.360 161.070 ;
        RECT 240.280 160.705 253.130 161.040 ;
        RECT 257.295 161.035 257.675 161.080 ;
        RECT 256.560 160.735 257.870 161.035 ;
        RECT 257.295 160.700 257.675 160.735 ;
        RECT 274.385 160.645 275.475 161.025 ;
        RECT 276.430 160.655 277.950 161.015 ;
        RECT 278.870 160.650 291.720 160.985 ;
        RECT 295.885 160.980 296.265 161.025 ;
        RECT 295.150 160.680 296.460 160.980 ;
        RECT 295.885 160.645 296.265 160.680 ;
        RECT 232.650 160.150 265.730 160.190 ;
        RECT 232.650 159.840 297.895 160.150 ;
        RECT 264.945 159.785 297.895 159.840 ;
        RECT 299.690 159.775 303.950 160.130 ;
        RECT 216.760 159.245 220.855 159.250 ;
        RECT 200.180 159.240 205.395 159.245 ;
        RECT 215.640 159.240 220.855 159.245 ;
        RECT 231.100 159.240 271.350 159.245 ;
        RECT 200.180 159.190 271.350 159.240 ;
        RECT 297.895 159.190 303.540 159.195 ;
        RECT 314.155 159.190 314.535 165.020 ;
        RECT 323.035 164.970 327.535 165.280 ;
        RECT 399.325 165.025 403.455 165.325 ;
        RECT 318.995 164.420 325.385 164.710 ;
        RECT 383.285 164.025 389.200 164.360 ;
        RECT 386.555 164.005 389.200 164.025 ;
        RECT 317.760 163.255 320.680 163.555 ;
        RECT 324.225 163.240 327.595 163.540 ;
        RECT 363.880 163.385 367.180 163.765 ;
        RECT 367.880 163.385 371.180 163.765 ;
        RECT 377.380 163.385 380.680 163.765 ;
        RECT 381.380 163.385 384.680 163.765 ;
        RECT 315.975 162.505 316.355 162.885 ;
        RECT 321.635 162.610 322.825 162.895 ;
        RECT 320.855 161.945 321.235 162.325 ;
        RECT 324.975 161.780 328.155 162.100 ;
        RECT 363.880 161.385 365.165 161.765 ;
        RECT 383.195 161.385 384.680 161.765 ;
        RECT 315.255 160.695 319.405 160.965 ;
        RECT 365.385 160.705 366.905 161.065 ;
        RECT 314.905 159.190 319.000 159.195 ;
        RECT 200.180 159.185 303.540 159.190 ;
        RECT 313.785 159.185 319.000 159.190 ;
        RECT 200.180 158.345 328.815 159.185 ;
        RECT 74.875 158.290 132.450 158.345 ;
        RECT 271.240 158.290 328.815 158.345 ;
        RECT 360.195 158.340 386.850 159.240 ;
        RECT 396.950 159.195 397.330 165.025 ;
        RECT 405.830 164.975 410.330 165.285 ;
        RECT 414.785 165.025 418.915 165.325 ;
        RECT 401.790 164.425 408.180 164.715 ;
        RECT 401.205 163.845 411.860 164.180 ;
        RECT 400.555 163.260 403.475 163.560 ;
        RECT 407.020 163.245 410.390 163.545 ;
        RECT 398.770 162.510 399.150 162.890 ;
        RECT 401.175 162.525 402.955 162.815 ;
        RECT 404.430 162.615 405.620 162.900 ;
        RECT 408.550 162.495 409.860 162.815 ;
        RECT 399.905 161.910 400.285 162.290 ;
        RECT 403.650 161.950 404.030 162.330 ;
        RECT 406.360 161.940 406.740 162.320 ;
        RECT 407.770 161.785 410.950 162.105 ;
        RECT 397.700 159.195 401.795 159.200 ;
        RECT 412.410 159.195 412.790 165.025 ;
        RECT 421.290 164.975 425.790 165.285 ;
        RECT 512.930 164.970 517.060 165.270 ;
        RECT 428.520 164.760 464.430 164.815 ;
        RECT 417.250 164.425 423.640 164.715 ;
        RECT 428.520 164.545 495.715 164.760 ;
        RECT 463.970 164.490 495.715 164.545 ;
        RECT 499.935 164.370 506.325 164.660 ;
        RECT 416.665 163.845 427.170 164.180 ;
        RECT 452.140 163.980 462.690 164.315 ;
        RECT 499.350 163.790 509.830 164.125 ;
        RECT 416.015 163.260 418.935 163.560 ;
        RECT 422.480 163.245 425.850 163.545 ;
        RECT 430.730 163.340 432.035 163.720 ;
        RECT 432.735 163.340 436.035 163.720 ;
        RECT 436.735 163.340 440.035 163.720 ;
        RECT 440.735 163.340 442.095 163.720 ;
        RECT 444.070 163.340 445.535 163.720 ;
        RECT 446.235 163.340 449.535 163.720 ;
        RECT 450.235 163.340 453.535 163.720 ;
        RECT 454.235 163.340 455.415 163.720 ;
        RECT 469.320 163.285 470.625 163.665 ;
        RECT 475.325 163.285 478.625 163.665 ;
        RECT 479.325 163.285 480.685 163.665 ;
        RECT 482.660 163.285 484.125 163.665 ;
        RECT 484.825 163.285 488.125 163.665 ;
        RECT 492.825 163.285 494.005 163.665 ;
        RECT 432.195 162.995 432.575 163.030 ;
        RECT 414.230 162.510 414.610 162.890 ;
        RECT 416.635 162.525 418.415 162.815 ;
        RECT 419.890 162.615 421.080 162.900 ;
        RECT 424.010 162.495 425.320 162.815 ;
        RECT 431.930 162.685 434.940 162.995 ;
        RECT 432.195 162.650 432.575 162.685 ;
        RECT 436.195 162.650 437.285 163.030 ;
        RECT 440.195 163.025 440.575 163.030 ;
        RECT 437.715 162.660 440.580 163.025 ;
        RECT 445.695 163.005 446.075 163.030 ;
        RECT 445.680 162.685 447.825 163.005 ;
        RECT 440.195 162.650 440.575 162.660 ;
        RECT 445.695 162.650 446.075 162.685 ;
        RECT 448.740 162.650 450.075 163.030 ;
        RECT 453.695 163.010 454.075 163.030 ;
        RECT 451.230 162.690 454.140 163.010 ;
        RECT 470.785 162.940 471.165 162.975 ;
        RECT 453.695 162.650 454.075 162.690 ;
        RECT 470.520 162.630 473.530 162.940 ;
        RECT 470.785 162.595 471.165 162.630 ;
        RECT 474.785 162.595 475.875 162.975 ;
        RECT 478.785 162.970 479.165 162.975 ;
        RECT 476.305 162.605 479.170 162.970 ;
        RECT 484.285 162.950 484.665 162.975 ;
        RECT 484.270 162.630 486.415 162.950 ;
        RECT 478.785 162.595 479.165 162.605 ;
        RECT 484.285 162.595 484.665 162.630 ;
        RECT 487.330 162.595 488.665 162.975 ;
        RECT 492.285 162.955 492.665 162.975 ;
        RECT 489.820 162.635 492.730 162.955 ;
        RECT 492.285 162.595 492.665 162.635 ;
        RECT 496.915 162.455 497.295 162.835 ;
        RECT 499.320 162.470 501.100 162.760 ;
        RECT 502.575 162.560 503.765 162.845 ;
        RECT 506.695 162.440 508.005 162.760 ;
        RECT 415.365 161.910 415.745 162.290 ;
        RECT 419.110 161.950 419.490 162.330 ;
        RECT 421.820 161.940 422.200 162.320 ;
        RECT 423.230 161.785 426.410 162.105 ;
        RECT 498.050 161.855 498.430 162.235 ;
        RECT 501.795 161.895 502.175 162.275 ;
        RECT 504.505 161.885 504.885 162.265 ;
        RECT 505.915 161.730 509.095 162.050 ;
        RECT 430.545 161.340 432.035 161.720 ;
        RECT 432.735 161.340 434.020 161.720 ;
        RECT 452.050 161.340 453.535 161.720 ;
        RECT 454.235 161.340 455.310 161.720 ;
        RECT 469.135 161.285 470.625 161.665 ;
        RECT 492.825 161.285 493.900 161.665 ;
        RECT 432.195 160.650 433.285 161.030 ;
        RECT 434.240 160.660 435.760 161.020 ;
        RECT 436.680 160.655 449.530 160.990 ;
        RECT 453.695 160.985 454.075 161.030 ;
        RECT 452.960 160.685 454.270 160.985 ;
        RECT 453.695 160.650 454.075 160.685 ;
        RECT 470.785 160.595 471.875 160.975 ;
        RECT 472.830 160.605 474.350 160.965 ;
        RECT 475.270 160.600 488.120 160.935 ;
        RECT 492.285 160.930 492.665 160.975 ;
        RECT 491.550 160.630 492.860 160.930 ;
        RECT 492.285 160.595 492.665 160.630 ;
        RECT 429.050 160.100 462.130 160.140 ;
        RECT 429.050 159.790 494.295 160.100 ;
        RECT 461.345 159.735 494.295 159.790 ;
        RECT 496.090 159.725 500.350 160.080 ;
        RECT 413.160 159.195 417.255 159.200 ;
        RECT 396.580 159.190 401.795 159.195 ;
        RECT 412.040 159.190 417.255 159.195 ;
        RECT 427.500 159.190 467.750 159.195 ;
        RECT 396.580 159.140 467.750 159.190 ;
        RECT 494.295 159.140 499.940 159.145 ;
        RECT 510.555 159.140 510.935 164.970 ;
        RECT 519.435 164.920 523.935 165.230 ;
        RECT 595.700 165.060 599.830 165.360 ;
        RECT 515.395 164.370 521.785 164.660 ;
        RECT 579.605 164.070 585.520 164.405 ;
        RECT 582.875 164.050 585.520 164.070 ;
        RECT 514.160 163.205 517.080 163.505 ;
        RECT 520.625 163.190 523.995 163.490 ;
        RECT 560.200 163.430 563.500 163.810 ;
        RECT 564.200 163.430 567.500 163.810 ;
        RECT 573.700 163.430 577.000 163.810 ;
        RECT 577.700 163.430 581.000 163.810 ;
        RECT 512.375 162.455 512.755 162.835 ;
        RECT 518.035 162.560 519.225 162.845 ;
        RECT 517.255 161.895 517.635 162.275 ;
        RECT 521.375 161.730 524.555 162.050 ;
        RECT 560.200 161.430 561.485 161.810 ;
        RECT 579.515 161.430 581.000 161.810 ;
        RECT 511.655 160.645 515.805 160.915 ;
        RECT 561.705 160.750 563.225 161.110 ;
        RECT 511.305 159.140 515.400 159.145 ;
        RECT 396.580 159.135 499.940 159.140 ;
        RECT 510.185 159.135 515.400 159.140 ;
        RECT 396.580 158.295 525.215 159.135 ;
        RECT 556.515 158.385 583.170 159.285 ;
        RECT 593.325 159.230 593.705 165.060 ;
        RECT 602.205 165.010 606.705 165.320 ;
        RECT 611.160 165.060 615.290 165.360 ;
        RECT 598.165 164.460 604.555 164.750 ;
        RECT 597.580 163.880 608.235 164.215 ;
        RECT 596.930 163.295 599.850 163.595 ;
        RECT 603.395 163.280 606.765 163.580 ;
        RECT 595.145 162.545 595.525 162.925 ;
        RECT 597.550 162.560 599.330 162.850 ;
        RECT 600.805 162.650 601.995 162.935 ;
        RECT 604.925 162.530 606.235 162.850 ;
        RECT 596.280 161.945 596.660 162.325 ;
        RECT 600.025 161.985 600.405 162.365 ;
        RECT 602.735 161.975 603.115 162.355 ;
        RECT 604.145 161.820 607.325 162.140 ;
        RECT 594.075 159.230 598.170 159.235 ;
        RECT 608.785 159.230 609.165 165.060 ;
        RECT 617.665 165.010 622.165 165.320 ;
        RECT 709.305 165.005 713.435 165.305 ;
        RECT 624.895 164.795 660.805 164.850 ;
        RECT 613.625 164.460 620.015 164.750 ;
        RECT 624.895 164.580 692.090 164.795 ;
        RECT 660.345 164.525 692.090 164.580 ;
        RECT 696.310 164.405 702.700 164.695 ;
        RECT 613.040 163.880 623.545 164.215 ;
        RECT 648.515 164.015 659.065 164.350 ;
        RECT 695.725 163.825 706.205 164.160 ;
        RECT 612.390 163.295 615.310 163.595 ;
        RECT 618.855 163.280 622.225 163.580 ;
        RECT 627.105 163.375 628.410 163.755 ;
        RECT 629.110 163.375 632.410 163.755 ;
        RECT 633.110 163.375 636.410 163.755 ;
        RECT 637.110 163.375 638.470 163.755 ;
        RECT 640.445 163.375 641.910 163.755 ;
        RECT 642.610 163.375 645.910 163.755 ;
        RECT 646.610 163.375 649.910 163.755 ;
        RECT 650.610 163.375 651.790 163.755 ;
        RECT 665.695 163.320 667.000 163.700 ;
        RECT 671.700 163.320 675.000 163.700 ;
        RECT 675.700 163.320 677.060 163.700 ;
        RECT 679.035 163.320 680.500 163.700 ;
        RECT 681.200 163.320 684.500 163.700 ;
        RECT 689.200 163.320 690.380 163.700 ;
        RECT 628.570 163.030 628.950 163.065 ;
        RECT 610.605 162.545 610.985 162.925 ;
        RECT 613.010 162.560 614.790 162.850 ;
        RECT 616.265 162.650 617.455 162.935 ;
        RECT 620.385 162.530 621.695 162.850 ;
        RECT 628.305 162.720 631.315 163.030 ;
        RECT 628.570 162.685 628.950 162.720 ;
        RECT 632.570 162.685 633.660 163.065 ;
        RECT 636.570 163.060 636.950 163.065 ;
        RECT 634.090 162.695 636.955 163.060 ;
        RECT 642.070 163.040 642.450 163.065 ;
        RECT 642.055 162.720 644.200 163.040 ;
        RECT 636.570 162.685 636.950 162.695 ;
        RECT 642.070 162.685 642.450 162.720 ;
        RECT 645.115 162.685 646.450 163.065 ;
        RECT 650.070 163.045 650.450 163.065 ;
        RECT 647.605 162.725 650.515 163.045 ;
        RECT 667.160 162.975 667.540 163.010 ;
        RECT 650.070 162.685 650.450 162.725 ;
        RECT 666.895 162.665 669.905 162.975 ;
        RECT 667.160 162.630 667.540 162.665 ;
        RECT 671.160 162.630 672.250 163.010 ;
        RECT 675.160 163.005 675.540 163.010 ;
        RECT 672.680 162.640 675.545 163.005 ;
        RECT 680.660 162.985 681.040 163.010 ;
        RECT 680.645 162.665 682.790 162.985 ;
        RECT 675.160 162.630 675.540 162.640 ;
        RECT 680.660 162.630 681.040 162.665 ;
        RECT 683.705 162.630 685.040 163.010 ;
        RECT 688.660 162.990 689.040 163.010 ;
        RECT 686.195 162.670 689.105 162.990 ;
        RECT 688.660 162.630 689.040 162.670 ;
        RECT 693.290 162.490 693.670 162.870 ;
        RECT 695.695 162.505 697.475 162.795 ;
        RECT 698.950 162.595 700.140 162.880 ;
        RECT 703.070 162.475 704.380 162.795 ;
        RECT 611.740 161.945 612.120 162.325 ;
        RECT 615.485 161.985 615.865 162.365 ;
        RECT 618.195 161.975 618.575 162.355 ;
        RECT 619.605 161.820 622.785 162.140 ;
        RECT 694.425 161.890 694.805 162.270 ;
        RECT 698.170 161.930 698.550 162.310 ;
        RECT 700.880 161.920 701.260 162.300 ;
        RECT 702.290 161.765 705.470 162.085 ;
        RECT 626.920 161.375 628.410 161.755 ;
        RECT 629.110 161.375 630.395 161.755 ;
        RECT 648.425 161.375 649.910 161.755 ;
        RECT 650.610 161.375 651.685 161.755 ;
        RECT 665.510 161.320 667.000 161.700 ;
        RECT 689.200 161.320 690.275 161.700 ;
        RECT 628.570 160.685 629.660 161.065 ;
        RECT 630.615 160.695 632.135 161.055 ;
        RECT 633.055 160.690 645.905 161.025 ;
        RECT 650.070 161.020 650.450 161.065 ;
        RECT 649.335 160.720 650.645 161.020 ;
        RECT 650.070 160.685 650.450 160.720 ;
        RECT 667.160 160.630 668.250 161.010 ;
        RECT 669.205 160.640 670.725 161.000 ;
        RECT 671.645 160.635 684.495 160.970 ;
        RECT 688.660 160.965 689.040 161.010 ;
        RECT 687.925 160.665 689.235 160.965 ;
        RECT 688.660 160.630 689.040 160.665 ;
        RECT 625.425 160.135 658.505 160.175 ;
        RECT 625.425 159.825 690.670 160.135 ;
        RECT 657.720 159.770 690.670 159.825 ;
        RECT 692.465 159.760 696.725 160.115 ;
        RECT 609.535 159.230 613.630 159.235 ;
        RECT 592.955 159.225 598.170 159.230 ;
        RECT 608.415 159.225 613.630 159.230 ;
        RECT 623.875 159.225 664.125 159.230 ;
        RECT 592.955 159.175 664.125 159.225 ;
        RECT 690.670 159.175 696.315 159.180 ;
        RECT 706.930 159.175 707.310 165.005 ;
        RECT 715.810 164.955 720.310 165.265 ;
        RECT 792.040 165.060 796.170 165.360 ;
        RECT 711.770 164.405 718.160 164.695 ;
        RECT 775.970 164.075 781.885 164.410 ;
        RECT 779.240 164.055 781.885 164.075 ;
        RECT 710.535 163.240 713.455 163.540 ;
        RECT 717.000 163.225 720.370 163.525 ;
        RECT 756.565 163.435 759.865 163.815 ;
        RECT 760.565 163.435 763.865 163.815 ;
        RECT 770.065 163.435 773.365 163.815 ;
        RECT 774.065 163.435 777.365 163.815 ;
        RECT 708.750 162.490 709.130 162.870 ;
        RECT 714.410 162.595 715.600 162.880 ;
        RECT 713.630 161.930 714.010 162.310 ;
        RECT 717.750 161.765 720.930 162.085 ;
        RECT 756.565 161.435 757.850 161.815 ;
        RECT 775.880 161.435 777.365 161.815 ;
        RECT 708.030 160.680 712.180 160.950 ;
        RECT 758.070 160.755 759.590 161.115 ;
        RECT 707.680 159.175 711.775 159.180 ;
        RECT 592.955 159.170 696.315 159.175 ;
        RECT 706.560 159.170 711.775 159.175 ;
        RECT 592.955 158.330 721.590 159.170 ;
        RECT 752.880 158.390 779.535 159.290 ;
        RECT 789.665 159.230 790.045 165.060 ;
        RECT 798.545 165.010 803.045 165.320 ;
        RECT 807.500 165.060 811.630 165.360 ;
        RECT 794.505 164.460 800.895 164.750 ;
        RECT 793.920 163.880 804.575 164.215 ;
        RECT 793.270 163.295 796.190 163.595 ;
        RECT 799.735 163.280 803.105 163.580 ;
        RECT 791.485 162.545 791.865 162.925 ;
        RECT 793.890 162.560 795.670 162.850 ;
        RECT 797.145 162.650 798.335 162.935 ;
        RECT 801.265 162.530 802.575 162.850 ;
        RECT 792.620 161.945 793.000 162.325 ;
        RECT 796.365 161.985 796.745 162.365 ;
        RECT 799.075 161.975 799.455 162.355 ;
        RECT 800.485 161.820 803.665 162.140 ;
        RECT 790.415 159.230 794.510 159.235 ;
        RECT 805.125 159.230 805.505 165.060 ;
        RECT 814.005 165.010 818.505 165.320 ;
        RECT 905.645 165.005 909.775 165.305 ;
        RECT 821.235 164.795 857.145 164.850 ;
        RECT 809.965 164.460 816.355 164.750 ;
        RECT 821.235 164.580 888.430 164.795 ;
        RECT 856.685 164.525 888.430 164.580 ;
        RECT 892.650 164.405 899.040 164.695 ;
        RECT 809.380 163.880 819.885 164.215 ;
        RECT 844.855 164.015 855.405 164.350 ;
        RECT 892.065 163.825 902.545 164.160 ;
        RECT 808.730 163.295 811.650 163.595 ;
        RECT 815.195 163.280 818.565 163.580 ;
        RECT 823.445 163.375 824.750 163.755 ;
        RECT 825.450 163.375 828.750 163.755 ;
        RECT 829.450 163.375 832.750 163.755 ;
        RECT 833.450 163.375 834.810 163.755 ;
        RECT 836.785 163.375 838.250 163.755 ;
        RECT 838.950 163.375 842.250 163.755 ;
        RECT 842.950 163.375 846.250 163.755 ;
        RECT 846.950 163.375 848.130 163.755 ;
        RECT 862.035 163.320 863.340 163.700 ;
        RECT 868.040 163.320 871.340 163.700 ;
        RECT 872.040 163.320 873.400 163.700 ;
        RECT 875.375 163.320 876.840 163.700 ;
        RECT 877.540 163.320 880.840 163.700 ;
        RECT 885.540 163.320 886.720 163.700 ;
        RECT 824.910 163.030 825.290 163.065 ;
        RECT 806.945 162.545 807.325 162.925 ;
        RECT 809.350 162.560 811.130 162.850 ;
        RECT 812.605 162.650 813.795 162.935 ;
        RECT 816.725 162.530 818.035 162.850 ;
        RECT 824.645 162.720 827.655 163.030 ;
        RECT 824.910 162.685 825.290 162.720 ;
        RECT 828.910 162.685 830.000 163.065 ;
        RECT 832.910 163.060 833.290 163.065 ;
        RECT 830.430 162.695 833.295 163.060 ;
        RECT 838.410 163.040 838.790 163.065 ;
        RECT 838.395 162.720 840.540 163.040 ;
        RECT 832.910 162.685 833.290 162.695 ;
        RECT 838.410 162.685 838.790 162.720 ;
        RECT 841.455 162.685 842.790 163.065 ;
        RECT 846.410 163.045 846.790 163.065 ;
        RECT 843.945 162.725 846.855 163.045 ;
        RECT 863.500 162.975 863.880 163.010 ;
        RECT 846.410 162.685 846.790 162.725 ;
        RECT 863.235 162.665 866.245 162.975 ;
        RECT 863.500 162.630 863.880 162.665 ;
        RECT 867.500 162.630 868.590 163.010 ;
        RECT 871.500 163.005 871.880 163.010 ;
        RECT 869.020 162.640 871.885 163.005 ;
        RECT 877.000 162.985 877.380 163.010 ;
        RECT 876.985 162.665 879.130 162.985 ;
        RECT 871.500 162.630 871.880 162.640 ;
        RECT 877.000 162.630 877.380 162.665 ;
        RECT 880.045 162.630 881.380 163.010 ;
        RECT 885.000 162.990 885.380 163.010 ;
        RECT 882.535 162.670 885.445 162.990 ;
        RECT 885.000 162.630 885.380 162.670 ;
        RECT 889.630 162.490 890.010 162.870 ;
        RECT 892.035 162.505 893.815 162.795 ;
        RECT 895.290 162.595 896.480 162.880 ;
        RECT 899.410 162.475 900.720 162.795 ;
        RECT 808.080 161.945 808.460 162.325 ;
        RECT 811.825 161.985 812.205 162.365 ;
        RECT 814.535 161.975 814.915 162.355 ;
        RECT 815.945 161.820 819.125 162.140 ;
        RECT 890.765 161.890 891.145 162.270 ;
        RECT 894.510 161.930 894.890 162.310 ;
        RECT 897.220 161.920 897.600 162.300 ;
        RECT 898.630 161.765 901.810 162.085 ;
        RECT 823.260 161.375 824.750 161.755 ;
        RECT 825.450 161.375 826.735 161.755 ;
        RECT 844.765 161.375 846.250 161.755 ;
        RECT 846.950 161.375 848.025 161.755 ;
        RECT 861.850 161.320 863.340 161.700 ;
        RECT 885.540 161.320 886.615 161.700 ;
        RECT 824.910 160.685 826.000 161.065 ;
        RECT 826.955 160.695 828.475 161.055 ;
        RECT 829.395 160.690 842.245 161.025 ;
        RECT 846.410 161.020 846.790 161.065 ;
        RECT 845.675 160.720 846.985 161.020 ;
        RECT 846.410 160.685 846.790 160.720 ;
        RECT 863.500 160.630 864.590 161.010 ;
        RECT 865.545 160.640 867.065 161.000 ;
        RECT 867.985 160.635 880.835 160.970 ;
        RECT 885.000 160.965 885.380 161.010 ;
        RECT 884.265 160.665 885.575 160.965 ;
        RECT 885.000 160.630 885.380 160.665 ;
        RECT 821.765 160.135 854.845 160.175 ;
        RECT 821.765 159.825 887.010 160.135 ;
        RECT 854.060 159.770 887.010 159.825 ;
        RECT 888.805 159.760 893.065 160.115 ;
        RECT 805.875 159.230 809.970 159.235 ;
        RECT 789.295 159.225 794.510 159.230 ;
        RECT 804.755 159.225 809.970 159.230 ;
        RECT 820.215 159.225 860.465 159.230 ;
        RECT 789.295 159.175 860.465 159.225 ;
        RECT 887.010 159.175 892.655 159.180 ;
        RECT 903.270 159.175 903.650 165.005 ;
        RECT 912.150 164.955 916.650 165.265 ;
        RECT 988.380 165.060 992.510 165.360 ;
        RECT 908.110 164.405 914.500 164.695 ;
        RECT 972.355 164.060 978.270 164.395 ;
        RECT 975.625 164.040 978.270 164.060 ;
        RECT 906.875 163.240 909.795 163.540 ;
        RECT 913.340 163.225 916.710 163.525 ;
        RECT 952.950 163.420 956.250 163.800 ;
        RECT 956.950 163.420 960.250 163.800 ;
        RECT 966.450 163.420 969.750 163.800 ;
        RECT 970.450 163.420 973.750 163.800 ;
        RECT 905.090 162.490 905.470 162.870 ;
        RECT 910.750 162.595 911.940 162.880 ;
        RECT 909.970 161.930 910.350 162.310 ;
        RECT 914.090 161.765 917.270 162.085 ;
        RECT 952.950 161.420 954.235 161.800 ;
        RECT 972.265 161.420 973.750 161.800 ;
        RECT 904.370 160.680 908.520 160.950 ;
        RECT 954.455 160.740 955.975 161.100 ;
        RECT 904.020 159.175 908.115 159.180 ;
        RECT 789.295 159.170 892.655 159.175 ;
        RECT 902.900 159.170 908.115 159.175 ;
        RECT 789.295 158.330 917.930 159.170 ;
        RECT 949.265 158.375 975.920 159.275 ;
        RECT 986.005 159.230 986.385 165.060 ;
        RECT 994.885 165.010 999.385 165.320 ;
        RECT 1003.840 165.060 1007.970 165.360 ;
        RECT 990.845 164.460 997.235 164.750 ;
        RECT 990.260 163.880 1000.915 164.215 ;
        RECT 989.610 163.295 992.530 163.595 ;
        RECT 996.075 163.280 999.445 163.580 ;
        RECT 987.825 162.545 988.205 162.925 ;
        RECT 990.230 162.560 992.010 162.850 ;
        RECT 993.485 162.650 994.675 162.935 ;
        RECT 997.605 162.530 998.915 162.850 ;
        RECT 988.960 161.945 989.340 162.325 ;
        RECT 992.705 161.985 993.085 162.365 ;
        RECT 995.415 161.975 995.795 162.355 ;
        RECT 996.825 161.820 1000.005 162.140 ;
        RECT 986.755 159.230 990.850 159.235 ;
        RECT 1001.465 159.230 1001.845 165.060 ;
        RECT 1010.345 165.010 1014.845 165.320 ;
        RECT 1101.985 165.005 1106.115 165.305 ;
        RECT 1017.575 164.795 1053.485 164.850 ;
        RECT 1006.305 164.460 1012.695 164.750 ;
        RECT 1017.575 164.580 1084.770 164.795 ;
        RECT 1053.025 164.525 1084.770 164.580 ;
        RECT 1088.990 164.405 1095.380 164.695 ;
        RECT 1005.720 163.880 1016.225 164.215 ;
        RECT 1041.195 164.015 1051.745 164.350 ;
        RECT 1088.405 163.825 1098.885 164.160 ;
        RECT 1005.070 163.295 1007.990 163.595 ;
        RECT 1011.535 163.280 1014.905 163.580 ;
        RECT 1019.785 163.375 1021.090 163.755 ;
        RECT 1021.790 163.375 1025.090 163.755 ;
        RECT 1025.790 163.375 1029.090 163.755 ;
        RECT 1029.790 163.375 1031.150 163.755 ;
        RECT 1033.125 163.375 1034.590 163.755 ;
        RECT 1035.290 163.375 1038.590 163.755 ;
        RECT 1039.290 163.375 1042.590 163.755 ;
        RECT 1043.290 163.375 1044.470 163.755 ;
        RECT 1058.375 163.320 1059.680 163.700 ;
        RECT 1064.380 163.320 1067.680 163.700 ;
        RECT 1068.380 163.320 1069.740 163.700 ;
        RECT 1071.715 163.320 1073.180 163.700 ;
        RECT 1073.880 163.320 1077.180 163.700 ;
        RECT 1081.880 163.320 1083.060 163.700 ;
        RECT 1021.250 163.030 1021.630 163.065 ;
        RECT 1003.285 162.545 1003.665 162.925 ;
        RECT 1005.690 162.560 1007.470 162.850 ;
        RECT 1008.945 162.650 1010.135 162.935 ;
        RECT 1013.065 162.530 1014.375 162.850 ;
        RECT 1020.985 162.720 1023.995 163.030 ;
        RECT 1021.250 162.685 1021.630 162.720 ;
        RECT 1025.250 162.685 1026.340 163.065 ;
        RECT 1029.250 163.060 1029.630 163.065 ;
        RECT 1026.770 162.695 1029.635 163.060 ;
        RECT 1034.750 163.040 1035.130 163.065 ;
        RECT 1034.735 162.720 1036.880 163.040 ;
        RECT 1029.250 162.685 1029.630 162.695 ;
        RECT 1034.750 162.685 1035.130 162.720 ;
        RECT 1037.795 162.685 1039.130 163.065 ;
        RECT 1042.750 163.045 1043.130 163.065 ;
        RECT 1040.285 162.725 1043.195 163.045 ;
        RECT 1059.840 162.975 1060.220 163.010 ;
        RECT 1042.750 162.685 1043.130 162.725 ;
        RECT 1059.575 162.665 1062.585 162.975 ;
        RECT 1059.840 162.630 1060.220 162.665 ;
        RECT 1063.840 162.630 1064.930 163.010 ;
        RECT 1067.840 163.005 1068.220 163.010 ;
        RECT 1065.360 162.640 1068.225 163.005 ;
        RECT 1073.340 162.985 1073.720 163.010 ;
        RECT 1073.325 162.665 1075.470 162.985 ;
        RECT 1067.840 162.630 1068.220 162.640 ;
        RECT 1073.340 162.630 1073.720 162.665 ;
        RECT 1076.385 162.630 1077.720 163.010 ;
        RECT 1081.340 162.990 1081.720 163.010 ;
        RECT 1078.875 162.670 1081.785 162.990 ;
        RECT 1081.340 162.630 1081.720 162.670 ;
        RECT 1085.970 162.490 1086.350 162.870 ;
        RECT 1088.375 162.505 1090.155 162.795 ;
        RECT 1091.630 162.595 1092.820 162.880 ;
        RECT 1095.750 162.475 1097.060 162.795 ;
        RECT 1004.420 161.945 1004.800 162.325 ;
        RECT 1008.165 161.985 1008.545 162.365 ;
        RECT 1010.875 161.975 1011.255 162.355 ;
        RECT 1012.285 161.820 1015.465 162.140 ;
        RECT 1087.105 161.890 1087.485 162.270 ;
        RECT 1090.850 161.930 1091.230 162.310 ;
        RECT 1093.560 161.920 1093.940 162.300 ;
        RECT 1094.970 161.765 1098.150 162.085 ;
        RECT 1019.600 161.375 1021.090 161.755 ;
        RECT 1021.790 161.375 1023.075 161.755 ;
        RECT 1041.105 161.375 1042.590 161.755 ;
        RECT 1043.290 161.375 1044.365 161.755 ;
        RECT 1058.190 161.320 1059.680 161.700 ;
        RECT 1081.880 161.320 1082.955 161.700 ;
        RECT 1021.250 160.685 1022.340 161.065 ;
        RECT 1023.295 160.695 1024.815 161.055 ;
        RECT 1025.735 160.690 1038.585 161.025 ;
        RECT 1042.750 161.020 1043.130 161.065 ;
        RECT 1042.015 160.720 1043.325 161.020 ;
        RECT 1042.750 160.685 1043.130 160.720 ;
        RECT 1059.840 160.630 1060.930 161.010 ;
        RECT 1061.885 160.640 1063.405 161.000 ;
        RECT 1064.325 160.635 1077.175 160.970 ;
        RECT 1081.340 160.965 1081.720 161.010 ;
        RECT 1080.605 160.665 1081.915 160.965 ;
        RECT 1081.340 160.630 1081.720 160.665 ;
        RECT 1018.105 160.135 1051.185 160.175 ;
        RECT 1018.105 159.825 1083.350 160.135 ;
        RECT 1050.400 159.770 1083.350 159.825 ;
        RECT 1085.145 159.760 1089.405 160.115 ;
        RECT 1002.215 159.230 1006.310 159.235 ;
        RECT 985.635 159.225 990.850 159.230 ;
        RECT 1001.095 159.225 1006.310 159.230 ;
        RECT 1016.555 159.225 1056.805 159.230 ;
        RECT 985.635 159.175 1056.805 159.225 ;
        RECT 1083.350 159.175 1088.995 159.180 ;
        RECT 1099.610 159.175 1099.990 165.005 ;
        RECT 1108.490 164.955 1112.990 165.265 ;
        RECT 1184.720 165.060 1188.850 165.360 ;
        RECT 1104.450 164.405 1110.840 164.695 ;
        RECT 1168.680 164.065 1174.595 164.400 ;
        RECT 1171.950 164.045 1174.595 164.065 ;
        RECT 1103.215 163.240 1106.135 163.540 ;
        RECT 1109.680 163.225 1113.050 163.525 ;
        RECT 1149.275 163.425 1152.575 163.805 ;
        RECT 1153.275 163.425 1156.575 163.805 ;
        RECT 1162.775 163.425 1166.075 163.805 ;
        RECT 1166.775 163.425 1170.075 163.805 ;
        RECT 1101.430 162.490 1101.810 162.870 ;
        RECT 1107.090 162.595 1108.280 162.880 ;
        RECT 1106.310 161.930 1106.690 162.310 ;
        RECT 1110.430 161.765 1113.610 162.085 ;
        RECT 1149.275 161.425 1150.560 161.805 ;
        RECT 1168.590 161.425 1170.075 161.805 ;
        RECT 1100.710 160.680 1104.860 160.950 ;
        RECT 1150.780 160.745 1152.300 161.105 ;
        RECT 1100.360 159.175 1104.455 159.180 ;
        RECT 985.635 159.170 1088.995 159.175 ;
        RECT 1099.240 159.170 1104.455 159.175 ;
        RECT 985.635 158.330 1114.270 159.170 ;
        RECT 1145.590 158.380 1172.245 159.280 ;
        RECT 1182.345 159.230 1182.725 165.060 ;
        RECT 1191.225 165.010 1195.725 165.320 ;
        RECT 1200.180 165.060 1204.310 165.360 ;
        RECT 1187.185 164.460 1193.575 164.750 ;
        RECT 1186.600 163.880 1197.255 164.215 ;
        RECT 1185.950 163.295 1188.870 163.595 ;
        RECT 1192.415 163.280 1195.785 163.580 ;
        RECT 1184.165 162.545 1184.545 162.925 ;
        RECT 1186.570 162.560 1188.350 162.850 ;
        RECT 1189.825 162.650 1191.015 162.935 ;
        RECT 1193.945 162.530 1195.255 162.850 ;
        RECT 1185.300 161.945 1185.680 162.325 ;
        RECT 1189.045 161.985 1189.425 162.365 ;
        RECT 1191.755 161.975 1192.135 162.355 ;
        RECT 1193.165 161.820 1196.345 162.140 ;
        RECT 1183.095 159.230 1187.190 159.235 ;
        RECT 1197.805 159.230 1198.185 165.060 ;
        RECT 1206.685 165.010 1211.185 165.320 ;
        RECT 1282.865 165.005 1286.995 165.305 ;
        RECT 1289.370 164.955 1293.870 165.265 ;
        RECT 1298.325 165.005 1302.455 165.305 ;
        RECT 1213.915 164.795 1249.825 164.850 ;
        RECT 1202.645 164.460 1209.035 164.750 ;
        RECT 1213.915 164.580 1281.110 164.795 ;
        RECT 1249.365 164.525 1281.110 164.580 ;
        RECT 1285.330 164.405 1291.720 164.695 ;
        RECT 1202.060 163.880 1212.565 164.215 ;
        RECT 1237.535 164.015 1248.085 164.350 ;
        RECT 1276.125 163.960 1280.070 164.295 ;
        RECT 1284.745 163.825 1295.225 164.160 ;
        RECT 1201.410 163.295 1204.330 163.595 ;
        RECT 1207.875 163.280 1211.245 163.580 ;
        RECT 1216.125 163.375 1217.430 163.755 ;
        RECT 1218.130 163.375 1221.430 163.755 ;
        RECT 1222.130 163.375 1225.430 163.755 ;
        RECT 1226.130 163.375 1227.490 163.755 ;
        RECT 1229.465 163.375 1230.930 163.755 ;
        RECT 1231.630 163.375 1234.930 163.755 ;
        RECT 1235.630 163.375 1238.930 163.755 ;
        RECT 1239.630 163.375 1240.810 163.755 ;
        RECT 1254.715 163.320 1256.020 163.700 ;
        RECT 1256.720 163.320 1260.020 163.700 ;
        RECT 1260.720 163.320 1264.020 163.700 ;
        RECT 1264.720 163.320 1266.080 163.700 ;
        RECT 1268.055 163.320 1269.520 163.700 ;
        RECT 1270.220 163.320 1273.520 163.700 ;
        RECT 1274.220 163.320 1277.520 163.700 ;
        RECT 1278.220 163.320 1279.400 163.700 ;
        RECT 1284.095 163.240 1287.015 163.540 ;
        RECT 1290.560 163.225 1293.930 163.525 ;
        RECT 1217.590 163.030 1217.970 163.065 ;
        RECT 1199.625 162.545 1200.005 162.925 ;
        RECT 1202.030 162.560 1203.810 162.850 ;
        RECT 1205.285 162.650 1206.475 162.935 ;
        RECT 1209.405 162.530 1210.715 162.850 ;
        RECT 1217.325 162.720 1220.335 163.030 ;
        RECT 1217.590 162.685 1217.970 162.720 ;
        RECT 1221.590 162.685 1222.680 163.065 ;
        RECT 1225.590 163.060 1225.970 163.065 ;
        RECT 1223.110 162.695 1225.975 163.060 ;
        RECT 1231.090 163.040 1231.470 163.065 ;
        RECT 1231.075 162.720 1233.220 163.040 ;
        RECT 1225.590 162.685 1225.970 162.695 ;
        RECT 1231.090 162.685 1231.470 162.720 ;
        RECT 1234.135 162.685 1235.470 163.065 ;
        RECT 1239.090 163.045 1239.470 163.065 ;
        RECT 1236.625 162.725 1239.535 163.045 ;
        RECT 1256.180 162.975 1256.560 163.010 ;
        RECT 1239.090 162.685 1239.470 162.725 ;
        RECT 1255.915 162.665 1258.925 162.975 ;
        RECT 1256.180 162.630 1256.560 162.665 ;
        RECT 1260.180 162.630 1261.270 163.010 ;
        RECT 1264.180 163.005 1264.560 163.010 ;
        RECT 1261.700 162.640 1264.565 163.005 ;
        RECT 1269.680 162.985 1270.060 163.010 ;
        RECT 1269.665 162.665 1271.810 162.985 ;
        RECT 1264.180 162.630 1264.560 162.640 ;
        RECT 1269.680 162.630 1270.060 162.665 ;
        RECT 1272.725 162.630 1274.060 163.010 ;
        RECT 1277.680 162.990 1278.060 163.010 ;
        RECT 1275.215 162.670 1278.125 162.990 ;
        RECT 1277.680 162.630 1278.060 162.670 ;
        RECT 1282.310 162.490 1282.690 162.870 ;
        RECT 1284.715 162.505 1286.495 162.795 ;
        RECT 1287.970 162.595 1289.160 162.880 ;
        RECT 1292.090 162.475 1293.400 162.795 ;
        RECT 1200.760 161.945 1201.140 162.325 ;
        RECT 1204.505 161.985 1204.885 162.365 ;
        RECT 1207.215 161.975 1207.595 162.355 ;
        RECT 1208.625 161.820 1211.805 162.140 ;
        RECT 1283.445 161.890 1283.825 162.270 ;
        RECT 1287.190 161.930 1287.570 162.310 ;
        RECT 1289.900 161.920 1290.280 162.300 ;
        RECT 1291.310 161.765 1294.490 162.085 ;
        RECT 1215.940 161.375 1217.430 161.755 ;
        RECT 1218.130 161.375 1219.415 161.755 ;
        RECT 1237.445 161.375 1238.930 161.755 ;
        RECT 1239.630 161.375 1240.705 161.755 ;
        RECT 1254.530 161.320 1256.020 161.700 ;
        RECT 1256.720 161.320 1258.005 161.700 ;
        RECT 1276.035 161.320 1277.520 161.700 ;
        RECT 1278.220 161.320 1279.295 161.700 ;
        RECT 1217.590 160.685 1218.680 161.065 ;
        RECT 1219.635 160.695 1221.155 161.055 ;
        RECT 1222.075 160.690 1234.925 161.025 ;
        RECT 1239.090 161.020 1239.470 161.065 ;
        RECT 1238.355 160.720 1239.665 161.020 ;
        RECT 1239.090 160.685 1239.470 160.720 ;
        RECT 1256.180 160.630 1257.270 161.010 ;
        RECT 1258.225 160.640 1259.745 161.000 ;
        RECT 1260.665 160.635 1273.515 160.970 ;
        RECT 1277.680 160.965 1278.060 161.010 ;
        RECT 1276.945 160.665 1278.255 160.965 ;
        RECT 1277.680 160.630 1278.060 160.665 ;
        RECT 1214.445 160.135 1247.525 160.175 ;
        RECT 1214.445 159.825 1279.690 160.135 ;
        RECT 1246.740 159.770 1279.690 159.825 ;
        RECT 1281.485 159.760 1285.745 160.115 ;
        RECT 1198.555 159.230 1202.650 159.235 ;
        RECT 1181.975 159.225 1187.190 159.230 ;
        RECT 1197.435 159.225 1202.650 159.230 ;
        RECT 1212.895 159.225 1253.145 159.230 ;
        RECT 1181.975 159.175 1253.145 159.225 ;
        RECT 1279.690 159.175 1285.335 159.180 ;
        RECT 1295.950 159.175 1296.330 165.005 ;
        RECT 1304.830 164.955 1309.330 165.265 ;
        RECT 1300.790 164.405 1307.180 164.695 ;
        RECT 1299.555 163.240 1302.475 163.540 ;
        RECT 1306.020 163.225 1309.390 163.525 ;
        RECT 1297.770 162.490 1298.150 162.870 ;
        RECT 1303.430 162.595 1304.620 162.880 ;
        RECT 1302.650 161.930 1303.030 162.310 ;
        RECT 1306.770 161.765 1309.950 162.085 ;
        RECT 1297.050 160.680 1301.200 160.950 ;
        RECT 1296.700 159.175 1300.795 159.180 ;
        RECT 1181.975 159.170 1285.335 159.175 ;
        RECT 1295.580 159.170 1300.795 159.175 ;
        RECT 1181.975 158.330 1310.610 159.170 ;
        RECT 467.640 158.240 525.215 158.295 ;
        RECT 664.015 158.275 721.590 158.330 ;
        RECT 860.355 158.275 917.930 158.330 ;
        RECT 1056.695 158.275 1114.270 158.330 ;
        RECT 1253.035 158.275 1310.610 158.330 ;
        RECT -81.555 153.600 -56.120 154.500 ;
        RECT -31.230 153.680 -5.795 154.580 ;
        RECT 3.770 154.490 76.160 154.580 ;
        RECT 3.770 153.680 132.250 154.490 ;
        RECT 164.940 153.690 190.375 154.590 ;
        RECT 200.135 154.490 272.525 154.580 ;
        RECT 200.135 153.680 328.615 154.490 ;
        RECT -79.070 151.420 -77.870 151.800 ;
        RECT -76.115 151.205 -73.840 151.715 ;
        RECT -71.215 151.205 -68.915 151.715 ;
        RECT -66.620 151.205 -64.340 151.715 ;
        RECT -59.545 151.520 -58.310 151.900 ;
        RECT -28.745 151.500 -27.545 151.880 ;
        RECT -25.790 151.285 -23.515 151.795 ;
        RECT -20.890 151.285 -18.590 151.795 ;
        RECT -16.295 151.285 -14.015 151.795 ;
        RECT -9.220 151.600 -7.985 151.980 ;
        RECT -79.070 149.120 -75.810 149.500 ;
        RECT -75.070 149.120 -71.810 149.500 ;
        RECT -65.570 149.120 -62.310 149.500 ;
        RECT -61.570 149.120 -58.310 149.500 ;
        RECT -28.745 149.200 -25.485 149.580 ;
        RECT -24.745 149.200 -21.485 149.580 ;
        RECT -15.245 149.200 -11.985 149.580 ;
        RECT -11.245 149.200 -7.985 149.580 ;
        RECT -78.405 147.535 -56.120 147.545 ;
        RECT -78.405 147.205 -54.580 147.535 ;
        RECT -28.080 147.285 -1.785 147.625 ;
        RECT -56.340 147.185 -54.580 147.205 ;
        RECT 4.140 146.520 4.520 153.680 ;
        RECT 5.970 149.465 9.345 149.865 ;
        RECT 9.715 149.225 10.095 149.605 ;
        RECT 12.430 149.265 12.810 149.645 ;
        RECT 16.615 149.215 16.995 149.595 ;
        RECT 7.040 148.800 8.780 149.090 ;
        RECT 10.830 148.750 12.030 149.040 ;
        RECT 13.540 148.720 16.150 149.145 ;
        RECT 17.750 148.815 18.130 149.195 ;
        RECT 5.285 148.040 18.850 148.355 ;
        RECT 5.280 147.295 18.840 147.595 ;
        RECT 5.300 146.580 12.025 146.880 ;
        RECT 15.725 146.280 18.830 146.555 ;
        RECT 19.600 146.520 19.980 153.680 ;
        RECT 75.895 153.590 132.250 153.680 ;
        RECT 36.240 152.605 73.790 152.695 ;
        RECT 36.240 152.410 101.655 152.605 ;
        RECT 72.880 152.320 101.655 152.410 ;
        RECT 103.325 152.300 110.030 152.600 ;
        RECT 37.750 151.500 39.205 151.880 ;
        RECT 39.945 151.500 41.145 151.880 ;
        RECT 42.900 151.285 45.175 151.795 ;
        RECT 47.800 151.285 50.100 151.795 ;
        RECT 52.395 151.285 54.675 151.795 ;
        RECT 59.470 151.600 60.705 151.980 ;
        RECT 61.445 151.600 62.725 151.980 ;
        RECT 76.185 151.410 77.640 151.790 ;
        RECT 60.885 151.245 61.265 151.280 ;
        RECT 39.385 151.140 39.765 151.180 ;
        RECT 39.315 150.835 42.150 151.140 ;
        RECT 58.130 150.935 61.265 151.245 ;
        RECT 81.335 151.195 83.610 151.705 ;
        RECT 86.235 151.195 88.535 151.705 ;
        RECT 90.830 151.195 93.110 151.705 ;
        RECT 99.880 151.510 101.160 151.890 ;
        RECT 99.320 151.155 99.700 151.190 ;
        RECT 77.820 151.050 78.200 151.090 ;
        RECT 60.885 150.900 61.265 150.935 ;
        RECT 39.385 150.800 39.765 150.835 ;
        RECT 77.750 150.745 80.585 151.050 ;
        RECT 96.565 150.845 99.700 151.155 ;
        RECT 99.320 150.810 99.700 150.845 ;
        RECT 77.820 150.710 78.200 150.745 ;
        RECT 21.430 149.425 24.835 149.865 ;
        RECT 25.175 149.225 25.555 149.605 ;
        RECT 27.890 149.265 28.270 149.645 ;
        RECT 32.075 149.215 32.455 149.595 ;
        RECT 37.910 149.200 39.205 149.580 ;
        RECT 39.945 149.200 43.205 149.580 ;
        RECT 43.945 149.200 47.205 149.580 ;
        RECT 47.945 149.200 49.130 149.580 ;
        RECT 51.395 149.200 52.705 149.580 ;
        RECT 53.445 149.200 56.705 149.580 ;
        RECT 57.445 149.200 60.705 149.580 ;
        RECT 61.445 149.200 62.460 149.580 ;
        RECT 22.500 148.800 24.240 149.090 ;
        RECT 26.290 148.750 27.490 149.040 ;
        RECT 29.000 148.720 31.595 149.095 ;
        RECT 33.210 148.815 33.590 149.195 ;
        RECT 76.345 149.110 77.640 149.490 ;
        RECT 82.380 149.110 85.640 149.490 ;
        RECT 86.380 149.110 87.565 149.490 ;
        RECT 89.830 149.110 91.140 149.490 ;
        RECT 91.880 149.110 95.140 149.490 ;
        RECT 99.880 149.110 100.895 149.490 ;
        RECT 103.960 149.355 107.375 149.775 ;
        RECT 107.705 149.135 108.085 149.515 ;
        RECT 110.420 149.175 110.800 149.555 ;
        RECT 114.605 149.125 114.985 149.505 ;
        RECT 39.385 148.500 39.765 148.880 ;
        RECT 43.385 148.500 43.765 148.880 ;
        RECT 47.385 148.835 47.765 148.880 ;
        RECT 52.885 148.835 53.265 148.880 ;
        RECT 47.335 148.520 53.270 148.835 ;
        RECT 47.385 148.500 47.765 148.520 ;
        RECT 52.885 148.500 53.265 148.520 ;
        RECT 56.885 148.500 57.265 148.880 ;
        RECT 60.885 148.500 61.265 148.880 ;
        RECT 77.820 148.410 78.200 148.790 ;
        RECT 81.820 148.410 82.200 148.790 ;
        RECT 85.820 148.745 86.200 148.790 ;
        RECT 91.320 148.745 91.700 148.790 ;
        RECT 85.770 148.430 91.705 148.745 ;
        RECT 85.820 148.410 86.200 148.430 ;
        RECT 91.320 148.410 91.700 148.430 ;
        RECT 95.320 148.410 95.700 148.790 ;
        RECT 99.320 148.410 99.700 148.790 ;
        RECT 105.030 148.710 106.770 149.000 ;
        RECT 108.820 148.660 110.020 148.950 ;
        RECT 111.530 148.620 114.160 149.075 ;
        RECT 115.740 148.725 116.120 149.105 ;
        RECT 20.740 148.040 34.565 148.340 ;
        RECT 36.240 147.875 52.250 148.250 ;
        RECT 69.910 147.785 90.685 148.160 ;
        RECT 20.745 147.295 39.165 147.595 ;
        RECT 40.610 147.285 67.920 147.625 ;
        RECT 20.225 146.580 27.485 146.880 ;
        RECT 5.280 145.960 9.405 146.230 ;
        RECT 20.780 146.045 24.865 146.315 ;
        RECT 31.185 146.280 34.935 146.555 ;
        RECT 36.240 146.520 62.470 146.910 ;
        RECT 68.940 146.430 100.905 146.820 ;
        RECT 113.715 146.190 116.845 146.465 ;
        RECT 117.590 146.430 117.970 153.590 ;
        RECT 167.425 151.510 168.625 151.890 ;
        RECT 118.830 151.130 125.570 151.430 ;
        RECT 170.380 151.295 172.655 151.805 ;
        RECT 175.280 151.295 177.580 151.805 ;
        RECT 179.875 151.295 182.155 151.805 ;
        RECT 186.950 151.610 188.185 151.990 ;
        RECT 119.420 149.335 122.875 149.775 ;
        RECT 123.165 149.135 123.545 149.515 ;
        RECT 125.880 149.175 126.260 149.555 ;
        RECT 130.065 149.125 130.445 149.505 ;
        RECT 167.425 149.210 170.685 149.590 ;
        RECT 171.425 149.210 174.685 149.590 ;
        RECT 180.925 149.210 184.185 149.590 ;
        RECT 184.925 149.210 188.185 149.590 ;
        RECT 120.490 148.710 122.230 149.000 ;
        RECT 124.280 148.660 125.480 148.950 ;
        RECT 126.990 148.630 129.615 149.040 ;
        RECT 131.200 148.725 131.580 149.105 ;
        RECT 118.235 147.950 134.155 148.250 ;
        RECT 118.770 147.205 135.715 147.505 ;
        RECT 168.090 147.295 194.385 147.635 ;
        RECT 200.505 146.520 200.885 153.680 ;
        RECT 202.335 149.465 205.710 149.865 ;
        RECT 206.080 149.225 206.460 149.605 ;
        RECT 208.795 149.265 209.175 149.645 ;
        RECT 212.980 149.215 213.360 149.595 ;
        RECT 203.405 148.800 205.145 149.090 ;
        RECT 207.195 148.750 208.395 149.040 ;
        RECT 209.905 148.720 212.515 149.145 ;
        RECT 214.115 148.815 214.495 149.195 ;
        RECT 201.650 148.040 215.215 148.355 ;
        RECT 201.645 147.295 215.205 147.595 ;
        RECT 201.665 146.580 208.390 146.880 ;
        RECT 129.175 146.190 136.875 146.465 ;
        RECT 212.090 146.280 215.195 146.555 ;
        RECT 215.965 146.520 216.345 153.680 ;
        RECT 272.260 153.590 328.615 153.680 ;
        RECT 361.330 153.650 386.765 154.550 ;
        RECT 396.535 154.440 468.925 154.530 ;
        RECT 396.535 153.630 525.015 154.440 ;
        RECT 557.650 153.695 583.085 154.595 ;
        RECT 592.910 154.475 665.300 154.565 ;
        RECT 592.910 153.665 721.390 154.475 ;
        RECT 754.015 153.700 779.450 154.600 ;
        RECT 789.250 154.475 861.640 154.565 ;
        RECT 789.250 153.665 917.730 154.475 ;
        RECT 950.400 153.685 975.835 154.585 ;
        RECT 985.590 154.475 1057.980 154.565 ;
        RECT 985.590 153.665 1114.070 154.475 ;
        RECT 1146.725 153.690 1172.160 154.590 ;
        RECT 1181.930 154.475 1254.320 154.565 ;
        RECT 1181.930 153.665 1310.410 154.475 ;
        RECT 232.605 152.605 270.155 152.695 ;
        RECT 232.605 152.410 298.020 152.605 ;
        RECT 269.245 152.320 298.020 152.410 ;
        RECT 299.690 152.300 306.395 152.600 ;
        RECT 234.115 151.500 235.570 151.880 ;
        RECT 236.310 151.500 237.510 151.880 ;
        RECT 239.265 151.285 241.540 151.795 ;
        RECT 244.165 151.285 246.465 151.795 ;
        RECT 248.760 151.285 251.040 151.795 ;
        RECT 255.835 151.600 257.070 151.980 ;
        RECT 257.810 151.600 259.090 151.980 ;
        RECT 272.550 151.410 274.005 151.790 ;
        RECT 257.250 151.245 257.630 151.280 ;
        RECT 235.750 151.140 236.130 151.180 ;
        RECT 235.680 150.835 238.515 151.140 ;
        RECT 254.495 150.935 257.630 151.245 ;
        RECT 277.700 151.195 279.975 151.705 ;
        RECT 282.600 151.195 284.900 151.705 ;
        RECT 287.195 151.195 289.475 151.705 ;
        RECT 296.245 151.510 297.525 151.890 ;
        RECT 295.685 151.155 296.065 151.190 ;
        RECT 274.185 151.050 274.565 151.090 ;
        RECT 257.250 150.900 257.630 150.935 ;
        RECT 235.750 150.800 236.130 150.835 ;
        RECT 274.115 150.745 276.950 151.050 ;
        RECT 292.930 150.845 296.065 151.155 ;
        RECT 295.685 150.810 296.065 150.845 ;
        RECT 274.185 150.710 274.565 150.745 ;
        RECT 217.795 149.425 221.200 149.865 ;
        RECT 221.540 149.225 221.920 149.605 ;
        RECT 224.255 149.265 224.635 149.645 ;
        RECT 228.440 149.215 228.820 149.595 ;
        RECT 234.275 149.200 235.570 149.580 ;
        RECT 236.310 149.200 239.570 149.580 ;
        RECT 240.310 149.200 243.570 149.580 ;
        RECT 244.310 149.200 245.495 149.580 ;
        RECT 247.760 149.200 249.070 149.580 ;
        RECT 249.810 149.200 253.070 149.580 ;
        RECT 253.810 149.200 257.070 149.580 ;
        RECT 257.810 149.200 258.825 149.580 ;
        RECT 218.865 148.800 220.605 149.090 ;
        RECT 222.655 148.750 223.855 149.040 ;
        RECT 225.365 148.720 227.960 149.095 ;
        RECT 229.575 148.815 229.955 149.195 ;
        RECT 272.710 149.110 274.005 149.490 ;
        RECT 278.745 149.110 282.005 149.490 ;
        RECT 282.745 149.110 283.930 149.490 ;
        RECT 286.195 149.110 287.505 149.490 ;
        RECT 288.245 149.110 291.505 149.490 ;
        RECT 296.245 149.110 297.260 149.490 ;
        RECT 300.325 149.355 303.740 149.775 ;
        RECT 304.070 149.135 304.450 149.515 ;
        RECT 306.785 149.175 307.165 149.555 ;
        RECT 310.970 149.125 311.350 149.505 ;
        RECT 235.750 148.500 236.130 148.880 ;
        RECT 239.750 148.500 240.130 148.880 ;
        RECT 243.750 148.835 244.130 148.880 ;
        RECT 249.250 148.835 249.630 148.880 ;
        RECT 243.700 148.520 249.635 148.835 ;
        RECT 243.750 148.500 244.130 148.520 ;
        RECT 249.250 148.500 249.630 148.520 ;
        RECT 253.250 148.500 253.630 148.880 ;
        RECT 257.250 148.500 257.630 148.880 ;
        RECT 274.185 148.410 274.565 148.790 ;
        RECT 278.185 148.410 278.565 148.790 ;
        RECT 282.185 148.745 282.565 148.790 ;
        RECT 287.685 148.745 288.065 148.790 ;
        RECT 282.135 148.430 288.070 148.745 ;
        RECT 282.185 148.410 282.565 148.430 ;
        RECT 287.685 148.410 288.065 148.430 ;
        RECT 291.685 148.410 292.065 148.790 ;
        RECT 295.685 148.410 296.065 148.790 ;
        RECT 301.395 148.710 303.135 149.000 ;
        RECT 305.185 148.660 306.385 148.950 ;
        RECT 307.895 148.620 310.525 149.075 ;
        RECT 312.105 148.725 312.485 149.105 ;
        RECT 217.105 148.040 230.930 148.340 ;
        RECT 232.605 147.875 248.615 148.250 ;
        RECT 266.275 147.785 287.050 148.160 ;
        RECT 217.110 147.295 235.530 147.595 ;
        RECT 236.975 147.285 264.285 147.625 ;
        RECT 216.590 146.580 223.850 146.880 ;
        RECT 36.240 146.155 54.910 146.165 ;
        RECT 36.240 146.075 66.260 146.155 ;
        RECT 36.240 146.065 93.345 146.075 ;
        RECT 36.240 145.845 102.350 146.065 ;
        RECT 201.645 145.960 205.770 146.230 ;
        RECT 217.145 146.045 221.230 146.315 ;
        RECT 227.550 146.280 231.300 146.555 ;
        RECT 232.605 146.520 258.835 146.910 ;
        RECT 265.305 146.430 297.270 146.820 ;
        RECT 310.080 146.190 313.210 146.465 ;
        RECT 313.955 146.430 314.335 153.590 ;
        RECT 363.815 151.470 365.015 151.850 ;
        RECT 315.195 151.130 321.935 151.430 ;
        RECT 366.770 151.255 369.045 151.765 ;
        RECT 371.670 151.255 373.970 151.765 ;
        RECT 376.265 151.255 378.545 151.765 ;
        RECT 383.340 151.570 384.575 151.950 ;
        RECT 315.785 149.335 319.240 149.775 ;
        RECT 319.530 149.135 319.910 149.515 ;
        RECT 322.245 149.175 322.625 149.555 ;
        RECT 326.430 149.125 326.810 149.505 ;
        RECT 363.815 149.170 367.075 149.550 ;
        RECT 367.815 149.170 371.075 149.550 ;
        RECT 377.315 149.170 380.575 149.550 ;
        RECT 381.315 149.170 384.575 149.550 ;
        RECT 316.855 148.710 318.595 149.000 ;
        RECT 320.645 148.660 321.845 148.950 ;
        RECT 323.355 148.630 325.980 149.040 ;
        RECT 327.565 148.725 327.945 149.105 ;
        RECT 314.600 147.950 330.520 148.250 ;
        RECT 315.135 147.205 332.080 147.505 ;
        RECT 364.480 147.255 390.775 147.595 ;
        RECT 396.905 146.470 397.285 153.630 ;
        RECT 398.735 149.415 402.110 149.815 ;
        RECT 402.480 149.175 402.860 149.555 ;
        RECT 405.195 149.215 405.575 149.595 ;
        RECT 409.380 149.165 409.760 149.545 ;
        RECT 399.805 148.750 401.545 149.040 ;
        RECT 403.595 148.700 404.795 148.990 ;
        RECT 406.305 148.670 408.915 149.095 ;
        RECT 410.515 148.765 410.895 149.145 ;
        RECT 398.050 147.990 411.615 148.305 ;
        RECT 398.045 147.245 411.605 147.545 ;
        RECT 398.065 146.530 404.790 146.830 ;
        RECT 325.540 146.190 333.240 146.465 ;
        RECT 408.490 146.230 411.595 146.505 ;
        RECT 412.365 146.470 412.745 153.630 ;
        RECT 468.660 153.540 525.015 153.630 ;
        RECT 429.005 152.555 466.555 152.645 ;
        RECT 429.005 152.360 494.420 152.555 ;
        RECT 465.645 152.270 494.420 152.360 ;
        RECT 496.090 152.250 502.795 152.550 ;
        RECT 430.515 151.450 431.970 151.830 ;
        RECT 432.710 151.450 433.910 151.830 ;
        RECT 435.665 151.235 437.940 151.745 ;
        RECT 440.565 151.235 442.865 151.745 ;
        RECT 445.160 151.235 447.440 151.745 ;
        RECT 452.235 151.550 453.470 151.930 ;
        RECT 454.210 151.550 455.490 151.930 ;
        RECT 468.950 151.360 470.405 151.740 ;
        RECT 453.650 151.195 454.030 151.230 ;
        RECT 432.150 151.090 432.530 151.130 ;
        RECT 432.080 150.785 434.915 151.090 ;
        RECT 450.895 150.885 454.030 151.195 ;
        RECT 474.100 151.145 476.375 151.655 ;
        RECT 479.000 151.145 481.300 151.655 ;
        RECT 483.595 151.145 485.875 151.655 ;
        RECT 492.645 151.460 493.925 151.840 ;
        RECT 492.085 151.105 492.465 151.140 ;
        RECT 470.585 151.000 470.965 151.040 ;
        RECT 453.650 150.850 454.030 150.885 ;
        RECT 432.150 150.750 432.530 150.785 ;
        RECT 470.515 150.695 473.350 151.000 ;
        RECT 489.330 150.795 492.465 151.105 ;
        RECT 492.085 150.760 492.465 150.795 ;
        RECT 470.585 150.660 470.965 150.695 ;
        RECT 414.195 149.375 417.600 149.815 ;
        RECT 417.940 149.175 418.320 149.555 ;
        RECT 420.655 149.215 421.035 149.595 ;
        RECT 424.840 149.165 425.220 149.545 ;
        RECT 430.675 149.150 431.970 149.530 ;
        RECT 432.710 149.150 435.970 149.530 ;
        RECT 436.710 149.150 439.970 149.530 ;
        RECT 440.710 149.150 441.895 149.530 ;
        RECT 444.160 149.150 445.470 149.530 ;
        RECT 446.210 149.150 449.470 149.530 ;
        RECT 450.210 149.150 453.470 149.530 ;
        RECT 454.210 149.150 455.225 149.530 ;
        RECT 415.265 148.750 417.005 149.040 ;
        RECT 419.055 148.700 420.255 148.990 ;
        RECT 421.765 148.670 424.360 149.045 ;
        RECT 425.975 148.765 426.355 149.145 ;
        RECT 469.110 149.060 470.405 149.440 ;
        RECT 475.145 149.060 478.405 149.440 ;
        RECT 479.145 149.060 480.330 149.440 ;
        RECT 482.595 149.060 483.905 149.440 ;
        RECT 484.645 149.060 487.905 149.440 ;
        RECT 492.645 149.060 493.660 149.440 ;
        RECT 496.725 149.305 500.140 149.725 ;
        RECT 500.470 149.085 500.850 149.465 ;
        RECT 503.185 149.125 503.565 149.505 ;
        RECT 507.370 149.075 507.750 149.455 ;
        RECT 432.150 148.450 432.530 148.830 ;
        RECT 436.150 148.450 436.530 148.830 ;
        RECT 440.150 148.785 440.530 148.830 ;
        RECT 445.650 148.785 446.030 148.830 ;
        RECT 440.100 148.470 446.035 148.785 ;
        RECT 440.150 148.450 440.530 148.470 ;
        RECT 445.650 148.450 446.030 148.470 ;
        RECT 449.650 148.450 450.030 148.830 ;
        RECT 453.650 148.450 454.030 148.830 ;
        RECT 470.585 148.360 470.965 148.740 ;
        RECT 474.585 148.360 474.965 148.740 ;
        RECT 478.585 148.695 478.965 148.740 ;
        RECT 484.085 148.695 484.465 148.740 ;
        RECT 478.535 148.380 484.470 148.695 ;
        RECT 478.585 148.360 478.965 148.380 ;
        RECT 484.085 148.360 484.465 148.380 ;
        RECT 488.085 148.360 488.465 148.740 ;
        RECT 492.085 148.360 492.465 148.740 ;
        RECT 497.795 148.660 499.535 148.950 ;
        RECT 501.585 148.610 502.785 148.900 ;
        RECT 504.295 148.570 506.925 149.025 ;
        RECT 508.505 148.675 508.885 149.055 ;
        RECT 413.505 147.990 427.330 148.290 ;
        RECT 429.005 147.825 445.015 148.200 ;
        RECT 462.675 147.735 483.450 148.110 ;
        RECT 413.510 147.245 431.930 147.545 ;
        RECT 433.375 147.235 460.685 147.575 ;
        RECT 412.990 146.530 420.250 146.830 ;
        RECT 232.605 146.155 251.275 146.165 ;
        RECT 232.605 146.075 262.625 146.155 ;
        RECT 232.605 146.065 289.710 146.075 ;
        RECT 232.605 145.845 298.715 146.065 ;
        RECT 398.045 145.910 402.170 146.180 ;
        RECT 413.545 145.995 417.630 146.265 ;
        RECT 423.950 146.230 427.700 146.505 ;
        RECT 429.005 146.470 455.235 146.860 ;
        RECT 461.705 146.380 493.670 146.770 ;
        RECT 506.480 146.140 509.610 146.415 ;
        RECT 510.355 146.380 510.735 153.540 ;
        RECT 560.135 151.515 561.335 151.895 ;
        RECT 511.595 151.080 518.335 151.380 ;
        RECT 563.090 151.300 565.365 151.810 ;
        RECT 567.990 151.300 570.290 151.810 ;
        RECT 572.585 151.300 574.865 151.810 ;
        RECT 579.660 151.615 580.895 151.995 ;
        RECT 512.185 149.285 515.640 149.725 ;
        RECT 515.930 149.085 516.310 149.465 ;
        RECT 518.645 149.125 519.025 149.505 ;
        RECT 522.830 149.075 523.210 149.455 ;
        RECT 560.135 149.215 563.395 149.595 ;
        RECT 564.135 149.215 567.395 149.595 ;
        RECT 573.635 149.215 576.895 149.595 ;
        RECT 577.635 149.215 580.895 149.595 ;
        RECT 513.255 148.660 514.995 148.950 ;
        RECT 517.045 148.610 518.245 148.900 ;
        RECT 519.755 148.580 522.380 148.990 ;
        RECT 523.965 148.675 524.345 149.055 ;
        RECT 511.000 147.900 526.920 148.200 ;
        RECT 511.535 147.155 528.480 147.455 ;
        RECT 560.800 147.300 587.095 147.640 ;
        RECT 593.280 146.505 593.660 153.665 ;
        RECT 595.110 149.450 598.485 149.850 ;
        RECT 598.855 149.210 599.235 149.590 ;
        RECT 601.570 149.250 601.950 149.630 ;
        RECT 605.755 149.200 606.135 149.580 ;
        RECT 596.180 148.785 597.920 149.075 ;
        RECT 599.970 148.735 601.170 149.025 ;
        RECT 602.680 148.705 605.290 149.130 ;
        RECT 606.890 148.800 607.270 149.180 ;
        RECT 594.425 148.025 607.990 148.340 ;
        RECT 594.420 147.280 607.980 147.580 ;
        RECT 594.440 146.565 601.165 146.865 ;
        RECT 521.940 146.140 529.640 146.415 ;
        RECT 604.865 146.265 607.970 146.540 ;
        RECT 608.740 146.505 609.120 153.665 ;
        RECT 665.035 153.575 721.390 153.665 ;
        RECT 625.380 152.590 662.930 152.680 ;
        RECT 625.380 152.395 690.795 152.590 ;
        RECT 662.020 152.305 690.795 152.395 ;
        RECT 692.465 152.285 699.170 152.585 ;
        RECT 626.890 151.485 628.345 151.865 ;
        RECT 629.085 151.485 630.285 151.865 ;
        RECT 632.040 151.270 634.315 151.780 ;
        RECT 636.940 151.270 639.240 151.780 ;
        RECT 641.535 151.270 643.815 151.780 ;
        RECT 648.610 151.585 649.845 151.965 ;
        RECT 650.585 151.585 651.865 151.965 ;
        RECT 665.325 151.395 666.780 151.775 ;
        RECT 650.025 151.230 650.405 151.265 ;
        RECT 628.525 151.125 628.905 151.165 ;
        RECT 628.455 150.820 631.290 151.125 ;
        RECT 647.270 150.920 650.405 151.230 ;
        RECT 670.475 151.180 672.750 151.690 ;
        RECT 675.375 151.180 677.675 151.690 ;
        RECT 679.970 151.180 682.250 151.690 ;
        RECT 689.020 151.495 690.300 151.875 ;
        RECT 688.460 151.140 688.840 151.175 ;
        RECT 666.960 151.035 667.340 151.075 ;
        RECT 650.025 150.885 650.405 150.920 ;
        RECT 628.525 150.785 628.905 150.820 ;
        RECT 666.890 150.730 669.725 151.035 ;
        RECT 685.705 150.830 688.840 151.140 ;
        RECT 688.460 150.795 688.840 150.830 ;
        RECT 666.960 150.695 667.340 150.730 ;
        RECT 610.570 149.410 613.975 149.850 ;
        RECT 614.315 149.210 614.695 149.590 ;
        RECT 617.030 149.250 617.410 149.630 ;
        RECT 621.215 149.200 621.595 149.580 ;
        RECT 627.050 149.185 628.345 149.565 ;
        RECT 629.085 149.185 632.345 149.565 ;
        RECT 633.085 149.185 636.345 149.565 ;
        RECT 637.085 149.185 638.270 149.565 ;
        RECT 640.535 149.185 641.845 149.565 ;
        RECT 642.585 149.185 645.845 149.565 ;
        RECT 646.585 149.185 649.845 149.565 ;
        RECT 650.585 149.185 651.600 149.565 ;
        RECT 611.640 148.785 613.380 149.075 ;
        RECT 615.430 148.735 616.630 149.025 ;
        RECT 618.140 148.705 620.735 149.080 ;
        RECT 622.350 148.800 622.730 149.180 ;
        RECT 665.485 149.095 666.780 149.475 ;
        RECT 671.520 149.095 674.780 149.475 ;
        RECT 675.520 149.095 676.705 149.475 ;
        RECT 678.970 149.095 680.280 149.475 ;
        RECT 681.020 149.095 684.280 149.475 ;
        RECT 689.020 149.095 690.035 149.475 ;
        RECT 693.100 149.340 696.515 149.760 ;
        RECT 696.845 149.120 697.225 149.500 ;
        RECT 699.560 149.160 699.940 149.540 ;
        RECT 703.745 149.110 704.125 149.490 ;
        RECT 628.525 148.485 628.905 148.865 ;
        RECT 632.525 148.485 632.905 148.865 ;
        RECT 636.525 148.820 636.905 148.865 ;
        RECT 642.025 148.820 642.405 148.865 ;
        RECT 636.475 148.505 642.410 148.820 ;
        RECT 636.525 148.485 636.905 148.505 ;
        RECT 642.025 148.485 642.405 148.505 ;
        RECT 646.025 148.485 646.405 148.865 ;
        RECT 650.025 148.485 650.405 148.865 ;
        RECT 666.960 148.395 667.340 148.775 ;
        RECT 670.960 148.395 671.340 148.775 ;
        RECT 674.960 148.730 675.340 148.775 ;
        RECT 680.460 148.730 680.840 148.775 ;
        RECT 674.910 148.415 680.845 148.730 ;
        RECT 674.960 148.395 675.340 148.415 ;
        RECT 680.460 148.395 680.840 148.415 ;
        RECT 684.460 148.395 684.840 148.775 ;
        RECT 688.460 148.395 688.840 148.775 ;
        RECT 694.170 148.695 695.910 148.985 ;
        RECT 697.960 148.645 699.160 148.935 ;
        RECT 700.670 148.605 703.300 149.060 ;
        RECT 704.880 148.710 705.260 149.090 ;
        RECT 609.880 148.025 623.705 148.325 ;
        RECT 625.380 147.860 641.390 148.235 ;
        RECT 659.050 147.770 679.825 148.145 ;
        RECT 609.885 147.280 628.305 147.580 ;
        RECT 629.750 147.270 657.060 147.610 ;
        RECT 609.365 146.565 616.625 146.865 ;
        RECT 429.005 146.105 447.675 146.115 ;
        RECT 429.005 146.025 459.025 146.105 ;
        RECT 429.005 146.015 486.110 146.025 ;
        RECT 65.785 145.755 102.350 145.845 ;
        RECT 262.150 145.755 298.715 145.845 ;
        RECT 429.005 145.795 495.115 146.015 ;
        RECT 594.420 145.945 598.545 146.215 ;
        RECT 609.920 146.030 614.005 146.300 ;
        RECT 620.325 146.265 624.075 146.540 ;
        RECT 625.380 146.505 651.610 146.895 ;
        RECT 658.080 146.415 690.045 146.805 ;
        RECT 702.855 146.175 705.985 146.450 ;
        RECT 706.730 146.415 707.110 153.575 ;
        RECT 756.500 151.520 757.700 151.900 ;
        RECT 707.970 151.115 714.710 151.415 ;
        RECT 759.455 151.305 761.730 151.815 ;
        RECT 764.355 151.305 766.655 151.815 ;
        RECT 768.950 151.305 771.230 151.815 ;
        RECT 776.025 151.620 777.260 152.000 ;
        RECT 708.560 149.320 712.015 149.760 ;
        RECT 712.305 149.120 712.685 149.500 ;
        RECT 715.020 149.160 715.400 149.540 ;
        RECT 719.205 149.110 719.585 149.490 ;
        RECT 756.500 149.220 759.760 149.600 ;
        RECT 760.500 149.220 763.760 149.600 ;
        RECT 770.000 149.220 773.260 149.600 ;
        RECT 774.000 149.220 777.260 149.600 ;
        RECT 709.630 148.695 711.370 148.985 ;
        RECT 713.420 148.645 714.620 148.935 ;
        RECT 716.130 148.615 718.755 149.025 ;
        RECT 720.340 148.710 720.720 149.090 ;
        RECT 707.375 147.935 723.295 148.235 ;
        RECT 707.910 147.190 724.855 147.490 ;
        RECT 757.165 147.305 783.460 147.645 ;
        RECT 789.620 146.505 790.000 153.665 ;
        RECT 791.450 149.450 794.825 149.850 ;
        RECT 795.195 149.210 795.575 149.590 ;
        RECT 797.910 149.250 798.290 149.630 ;
        RECT 802.095 149.200 802.475 149.580 ;
        RECT 792.520 148.785 794.260 149.075 ;
        RECT 796.310 148.735 797.510 149.025 ;
        RECT 799.020 148.705 801.630 149.130 ;
        RECT 803.230 148.800 803.610 149.180 ;
        RECT 790.765 148.025 804.330 148.340 ;
        RECT 790.760 147.280 804.320 147.580 ;
        RECT 790.780 146.565 797.505 146.865 ;
        RECT 718.315 146.175 726.015 146.450 ;
        RECT 801.205 146.265 804.310 146.540 ;
        RECT 805.080 146.505 805.460 153.665 ;
        RECT 861.375 153.575 917.730 153.665 ;
        RECT 821.720 152.590 859.270 152.680 ;
        RECT 821.720 152.395 887.135 152.590 ;
        RECT 858.360 152.305 887.135 152.395 ;
        RECT 888.805 152.285 895.510 152.585 ;
        RECT 823.230 151.485 824.685 151.865 ;
        RECT 825.425 151.485 826.625 151.865 ;
        RECT 828.380 151.270 830.655 151.780 ;
        RECT 833.280 151.270 835.580 151.780 ;
        RECT 837.875 151.270 840.155 151.780 ;
        RECT 844.950 151.585 846.185 151.965 ;
        RECT 846.925 151.585 848.205 151.965 ;
        RECT 861.665 151.395 863.120 151.775 ;
        RECT 846.365 151.230 846.745 151.265 ;
        RECT 824.865 151.125 825.245 151.165 ;
        RECT 824.795 150.820 827.630 151.125 ;
        RECT 843.610 150.920 846.745 151.230 ;
        RECT 866.815 151.180 869.090 151.690 ;
        RECT 871.715 151.180 874.015 151.690 ;
        RECT 876.310 151.180 878.590 151.690 ;
        RECT 885.360 151.495 886.640 151.875 ;
        RECT 884.800 151.140 885.180 151.175 ;
        RECT 863.300 151.035 863.680 151.075 ;
        RECT 846.365 150.885 846.745 150.920 ;
        RECT 824.865 150.785 825.245 150.820 ;
        RECT 863.230 150.730 866.065 151.035 ;
        RECT 882.045 150.830 885.180 151.140 ;
        RECT 884.800 150.795 885.180 150.830 ;
        RECT 863.300 150.695 863.680 150.730 ;
        RECT 806.910 149.410 810.315 149.850 ;
        RECT 810.655 149.210 811.035 149.590 ;
        RECT 813.370 149.250 813.750 149.630 ;
        RECT 817.555 149.200 817.935 149.580 ;
        RECT 823.390 149.185 824.685 149.565 ;
        RECT 825.425 149.185 828.685 149.565 ;
        RECT 829.425 149.185 832.685 149.565 ;
        RECT 833.425 149.185 834.610 149.565 ;
        RECT 836.875 149.185 838.185 149.565 ;
        RECT 838.925 149.185 842.185 149.565 ;
        RECT 842.925 149.185 846.185 149.565 ;
        RECT 846.925 149.185 847.940 149.565 ;
        RECT 807.980 148.785 809.720 149.075 ;
        RECT 811.770 148.735 812.970 149.025 ;
        RECT 814.480 148.705 817.075 149.080 ;
        RECT 818.690 148.800 819.070 149.180 ;
        RECT 861.825 149.095 863.120 149.475 ;
        RECT 867.860 149.095 871.120 149.475 ;
        RECT 871.860 149.095 873.045 149.475 ;
        RECT 875.310 149.095 876.620 149.475 ;
        RECT 877.360 149.095 880.620 149.475 ;
        RECT 885.360 149.095 886.375 149.475 ;
        RECT 889.440 149.340 892.855 149.760 ;
        RECT 893.185 149.120 893.565 149.500 ;
        RECT 895.900 149.160 896.280 149.540 ;
        RECT 900.085 149.110 900.465 149.490 ;
        RECT 824.865 148.485 825.245 148.865 ;
        RECT 828.865 148.485 829.245 148.865 ;
        RECT 832.865 148.820 833.245 148.865 ;
        RECT 838.365 148.820 838.745 148.865 ;
        RECT 832.815 148.505 838.750 148.820 ;
        RECT 832.865 148.485 833.245 148.505 ;
        RECT 838.365 148.485 838.745 148.505 ;
        RECT 842.365 148.485 842.745 148.865 ;
        RECT 846.365 148.485 846.745 148.865 ;
        RECT 863.300 148.395 863.680 148.775 ;
        RECT 867.300 148.395 867.680 148.775 ;
        RECT 871.300 148.730 871.680 148.775 ;
        RECT 876.800 148.730 877.180 148.775 ;
        RECT 871.250 148.415 877.185 148.730 ;
        RECT 871.300 148.395 871.680 148.415 ;
        RECT 876.800 148.395 877.180 148.415 ;
        RECT 880.800 148.395 881.180 148.775 ;
        RECT 884.800 148.395 885.180 148.775 ;
        RECT 890.510 148.695 892.250 148.985 ;
        RECT 894.300 148.645 895.500 148.935 ;
        RECT 897.010 148.605 899.640 149.060 ;
        RECT 901.220 148.710 901.600 149.090 ;
        RECT 806.220 148.025 820.045 148.325 ;
        RECT 821.720 147.860 837.730 148.235 ;
        RECT 855.390 147.770 876.165 148.145 ;
        RECT 806.225 147.280 824.645 147.580 ;
        RECT 826.090 147.270 853.400 147.610 ;
        RECT 805.705 146.565 812.965 146.865 ;
        RECT 625.380 146.140 644.050 146.150 ;
        RECT 625.380 146.060 655.400 146.140 ;
        RECT 625.380 146.050 682.485 146.060 ;
        RECT 625.380 145.830 691.490 146.050 ;
        RECT 790.760 145.945 794.885 146.215 ;
        RECT 806.260 146.030 810.345 146.300 ;
        RECT 816.665 146.265 820.415 146.540 ;
        RECT 821.720 146.505 847.950 146.895 ;
        RECT 854.420 146.415 886.385 146.805 ;
        RECT 899.195 146.175 902.325 146.450 ;
        RECT 903.070 146.415 903.450 153.575 ;
        RECT 952.885 151.505 954.085 151.885 ;
        RECT 904.310 151.115 911.050 151.415 ;
        RECT 955.840 151.290 958.115 151.800 ;
        RECT 960.740 151.290 963.040 151.800 ;
        RECT 965.335 151.290 967.615 151.800 ;
        RECT 972.410 151.605 973.645 151.985 ;
        RECT 904.900 149.320 908.355 149.760 ;
        RECT 908.645 149.120 909.025 149.500 ;
        RECT 911.360 149.160 911.740 149.540 ;
        RECT 915.545 149.110 915.925 149.490 ;
        RECT 952.885 149.205 956.145 149.585 ;
        RECT 956.885 149.205 960.145 149.585 ;
        RECT 966.385 149.205 969.645 149.585 ;
        RECT 970.385 149.205 973.645 149.585 ;
        RECT 905.970 148.695 907.710 148.985 ;
        RECT 909.760 148.645 910.960 148.935 ;
        RECT 912.470 148.615 915.095 149.025 ;
        RECT 916.680 148.710 917.060 149.090 ;
        RECT 903.715 147.935 919.635 148.235 ;
        RECT 904.250 147.190 921.195 147.490 ;
        RECT 953.550 147.290 979.845 147.630 ;
        RECT 985.960 146.505 986.340 153.665 ;
        RECT 987.790 149.450 991.165 149.850 ;
        RECT 991.535 149.210 991.915 149.590 ;
        RECT 994.250 149.250 994.630 149.630 ;
        RECT 998.435 149.200 998.815 149.580 ;
        RECT 988.860 148.785 990.600 149.075 ;
        RECT 992.650 148.735 993.850 149.025 ;
        RECT 995.360 148.705 997.970 149.130 ;
        RECT 999.570 148.800 999.950 149.180 ;
        RECT 987.105 148.025 1000.670 148.340 ;
        RECT 987.100 147.280 1000.660 147.580 ;
        RECT 987.120 146.565 993.845 146.865 ;
        RECT 914.655 146.175 922.355 146.450 ;
        RECT 997.545 146.265 1000.650 146.540 ;
        RECT 1001.420 146.505 1001.800 153.665 ;
        RECT 1057.715 153.575 1114.070 153.665 ;
        RECT 1018.060 152.590 1055.610 152.680 ;
        RECT 1018.060 152.395 1083.475 152.590 ;
        RECT 1054.700 152.305 1083.475 152.395 ;
        RECT 1085.145 152.285 1091.850 152.585 ;
        RECT 1019.570 151.485 1021.025 151.865 ;
        RECT 1021.765 151.485 1022.965 151.865 ;
        RECT 1024.720 151.270 1026.995 151.780 ;
        RECT 1029.620 151.270 1031.920 151.780 ;
        RECT 1034.215 151.270 1036.495 151.780 ;
        RECT 1041.290 151.585 1042.525 151.965 ;
        RECT 1043.265 151.585 1044.545 151.965 ;
        RECT 1058.005 151.395 1059.460 151.775 ;
        RECT 1042.705 151.230 1043.085 151.265 ;
        RECT 1021.205 151.125 1021.585 151.165 ;
        RECT 1021.135 150.820 1023.970 151.125 ;
        RECT 1039.950 150.920 1043.085 151.230 ;
        RECT 1063.155 151.180 1065.430 151.690 ;
        RECT 1068.055 151.180 1070.355 151.690 ;
        RECT 1072.650 151.180 1074.930 151.690 ;
        RECT 1081.700 151.495 1082.980 151.875 ;
        RECT 1081.140 151.140 1081.520 151.175 ;
        RECT 1059.640 151.035 1060.020 151.075 ;
        RECT 1042.705 150.885 1043.085 150.920 ;
        RECT 1021.205 150.785 1021.585 150.820 ;
        RECT 1059.570 150.730 1062.405 151.035 ;
        RECT 1078.385 150.830 1081.520 151.140 ;
        RECT 1081.140 150.795 1081.520 150.830 ;
        RECT 1059.640 150.695 1060.020 150.730 ;
        RECT 1003.250 149.410 1006.655 149.850 ;
        RECT 1006.995 149.210 1007.375 149.590 ;
        RECT 1009.710 149.250 1010.090 149.630 ;
        RECT 1013.895 149.200 1014.275 149.580 ;
        RECT 1019.730 149.185 1021.025 149.565 ;
        RECT 1021.765 149.185 1025.025 149.565 ;
        RECT 1025.765 149.185 1029.025 149.565 ;
        RECT 1029.765 149.185 1030.950 149.565 ;
        RECT 1033.215 149.185 1034.525 149.565 ;
        RECT 1035.265 149.185 1038.525 149.565 ;
        RECT 1039.265 149.185 1042.525 149.565 ;
        RECT 1043.265 149.185 1044.280 149.565 ;
        RECT 1004.320 148.785 1006.060 149.075 ;
        RECT 1008.110 148.735 1009.310 149.025 ;
        RECT 1010.820 148.705 1013.415 149.080 ;
        RECT 1015.030 148.800 1015.410 149.180 ;
        RECT 1058.165 149.095 1059.460 149.475 ;
        RECT 1064.200 149.095 1067.460 149.475 ;
        RECT 1068.200 149.095 1069.385 149.475 ;
        RECT 1071.650 149.095 1072.960 149.475 ;
        RECT 1073.700 149.095 1076.960 149.475 ;
        RECT 1081.700 149.095 1082.715 149.475 ;
        RECT 1085.780 149.340 1089.195 149.760 ;
        RECT 1089.525 149.120 1089.905 149.500 ;
        RECT 1092.240 149.160 1092.620 149.540 ;
        RECT 1096.425 149.110 1096.805 149.490 ;
        RECT 1021.205 148.485 1021.585 148.865 ;
        RECT 1025.205 148.485 1025.585 148.865 ;
        RECT 1029.205 148.820 1029.585 148.865 ;
        RECT 1034.705 148.820 1035.085 148.865 ;
        RECT 1029.155 148.505 1035.090 148.820 ;
        RECT 1029.205 148.485 1029.585 148.505 ;
        RECT 1034.705 148.485 1035.085 148.505 ;
        RECT 1038.705 148.485 1039.085 148.865 ;
        RECT 1042.705 148.485 1043.085 148.865 ;
        RECT 1059.640 148.395 1060.020 148.775 ;
        RECT 1063.640 148.395 1064.020 148.775 ;
        RECT 1067.640 148.730 1068.020 148.775 ;
        RECT 1073.140 148.730 1073.520 148.775 ;
        RECT 1067.590 148.415 1073.525 148.730 ;
        RECT 1067.640 148.395 1068.020 148.415 ;
        RECT 1073.140 148.395 1073.520 148.415 ;
        RECT 1077.140 148.395 1077.520 148.775 ;
        RECT 1081.140 148.395 1081.520 148.775 ;
        RECT 1086.850 148.695 1088.590 148.985 ;
        RECT 1090.640 148.645 1091.840 148.935 ;
        RECT 1093.350 148.605 1095.980 149.060 ;
        RECT 1097.560 148.710 1097.940 149.090 ;
        RECT 1002.560 148.025 1016.385 148.325 ;
        RECT 1018.060 147.860 1034.070 148.235 ;
        RECT 1051.730 147.770 1072.505 148.145 ;
        RECT 1002.565 147.280 1020.985 147.580 ;
        RECT 1022.430 147.270 1049.740 147.610 ;
        RECT 1002.045 146.565 1009.305 146.865 ;
        RECT 821.720 146.140 840.390 146.150 ;
        RECT 821.720 146.060 851.740 146.140 ;
        RECT 821.720 146.050 878.825 146.060 ;
        RECT 821.720 145.830 887.830 146.050 ;
        RECT 987.100 145.945 991.225 146.215 ;
        RECT 1002.600 146.030 1006.685 146.300 ;
        RECT 1013.005 146.265 1016.755 146.540 ;
        RECT 1018.060 146.505 1044.290 146.895 ;
        RECT 1050.760 146.415 1082.725 146.805 ;
        RECT 1095.535 146.175 1098.665 146.450 ;
        RECT 1099.410 146.415 1099.790 153.575 ;
        RECT 1149.210 151.510 1150.410 151.890 ;
        RECT 1100.650 151.115 1107.390 151.415 ;
        RECT 1152.165 151.295 1154.440 151.805 ;
        RECT 1157.065 151.295 1159.365 151.805 ;
        RECT 1161.660 151.295 1163.940 151.805 ;
        RECT 1168.735 151.610 1169.970 151.990 ;
        RECT 1101.240 149.320 1104.695 149.760 ;
        RECT 1104.985 149.120 1105.365 149.500 ;
        RECT 1107.700 149.160 1108.080 149.540 ;
        RECT 1111.885 149.110 1112.265 149.490 ;
        RECT 1149.210 149.210 1152.470 149.590 ;
        RECT 1153.210 149.210 1156.470 149.590 ;
        RECT 1162.710 149.210 1165.970 149.590 ;
        RECT 1166.710 149.210 1169.970 149.590 ;
        RECT 1102.310 148.695 1104.050 148.985 ;
        RECT 1106.100 148.645 1107.300 148.935 ;
        RECT 1108.810 148.615 1111.435 149.025 ;
        RECT 1113.020 148.710 1113.400 149.090 ;
        RECT 1100.055 147.935 1115.975 148.235 ;
        RECT 1100.590 147.190 1117.535 147.490 ;
        RECT 1149.875 147.295 1176.170 147.635 ;
        RECT 1182.300 146.505 1182.680 153.665 ;
        RECT 1184.130 149.450 1187.505 149.850 ;
        RECT 1187.875 149.210 1188.255 149.590 ;
        RECT 1190.590 149.250 1190.970 149.630 ;
        RECT 1194.775 149.200 1195.155 149.580 ;
        RECT 1185.200 148.785 1186.940 149.075 ;
        RECT 1188.990 148.735 1190.190 149.025 ;
        RECT 1191.700 148.705 1194.310 149.130 ;
        RECT 1195.910 148.800 1196.290 149.180 ;
        RECT 1183.445 148.025 1197.010 148.340 ;
        RECT 1183.440 147.280 1197.000 147.580 ;
        RECT 1183.460 146.565 1190.185 146.865 ;
        RECT 1110.995 146.175 1118.695 146.450 ;
        RECT 1193.885 146.265 1196.990 146.540 ;
        RECT 1197.760 146.505 1198.140 153.665 ;
        RECT 1254.055 153.575 1310.410 153.665 ;
        RECT 1214.400 152.590 1251.950 152.680 ;
        RECT 1214.400 152.395 1279.815 152.590 ;
        RECT 1251.040 152.305 1279.815 152.395 ;
        RECT 1281.485 152.285 1288.190 152.585 ;
        RECT 1215.910 151.485 1217.365 151.865 ;
        RECT 1218.105 151.485 1219.305 151.865 ;
        RECT 1221.060 151.270 1223.335 151.780 ;
        RECT 1225.960 151.270 1228.260 151.780 ;
        RECT 1230.555 151.270 1232.835 151.780 ;
        RECT 1237.630 151.585 1238.865 151.965 ;
        RECT 1239.605 151.585 1240.885 151.965 ;
        RECT 1254.345 151.395 1255.800 151.775 ;
        RECT 1256.540 151.395 1257.740 151.775 ;
        RECT 1239.045 151.230 1239.425 151.265 ;
        RECT 1217.545 151.125 1217.925 151.165 ;
        RECT 1217.475 150.820 1220.310 151.125 ;
        RECT 1236.290 150.920 1239.425 151.230 ;
        RECT 1259.495 151.180 1261.770 151.690 ;
        RECT 1264.395 151.180 1266.695 151.690 ;
        RECT 1268.990 151.180 1271.270 151.690 ;
        RECT 1276.065 151.495 1277.300 151.875 ;
        RECT 1278.040 151.495 1279.320 151.875 ;
        RECT 1277.480 151.140 1277.860 151.175 ;
        RECT 1255.980 151.035 1256.360 151.075 ;
        RECT 1239.045 150.885 1239.425 150.920 ;
        RECT 1217.545 150.785 1217.925 150.820 ;
        RECT 1255.910 150.730 1258.745 151.035 ;
        RECT 1274.725 150.830 1277.860 151.140 ;
        RECT 1277.480 150.795 1277.860 150.830 ;
        RECT 1255.980 150.695 1256.360 150.730 ;
        RECT 1199.590 149.410 1202.995 149.850 ;
        RECT 1203.335 149.210 1203.715 149.590 ;
        RECT 1206.050 149.250 1206.430 149.630 ;
        RECT 1210.235 149.200 1210.615 149.580 ;
        RECT 1216.070 149.185 1217.365 149.565 ;
        RECT 1218.105 149.185 1221.365 149.565 ;
        RECT 1222.105 149.185 1225.365 149.565 ;
        RECT 1226.105 149.185 1227.290 149.565 ;
        RECT 1229.555 149.185 1230.865 149.565 ;
        RECT 1231.605 149.185 1234.865 149.565 ;
        RECT 1235.605 149.185 1238.865 149.565 ;
        RECT 1239.605 149.185 1240.620 149.565 ;
        RECT 1200.660 148.785 1202.400 149.075 ;
        RECT 1204.450 148.735 1205.650 149.025 ;
        RECT 1207.160 148.705 1209.755 149.080 ;
        RECT 1211.370 148.800 1211.750 149.180 ;
        RECT 1254.505 149.095 1255.800 149.475 ;
        RECT 1256.540 149.095 1259.800 149.475 ;
        RECT 1260.540 149.095 1263.800 149.475 ;
        RECT 1264.540 149.095 1265.725 149.475 ;
        RECT 1267.990 149.095 1269.300 149.475 ;
        RECT 1270.040 149.095 1273.300 149.475 ;
        RECT 1274.040 149.095 1277.300 149.475 ;
        RECT 1278.040 149.095 1279.055 149.475 ;
        RECT 1282.120 149.340 1285.535 149.760 ;
        RECT 1285.865 149.120 1286.245 149.500 ;
        RECT 1288.580 149.160 1288.960 149.540 ;
        RECT 1292.765 149.110 1293.145 149.490 ;
        RECT 1217.545 148.485 1217.925 148.865 ;
        RECT 1221.545 148.485 1221.925 148.865 ;
        RECT 1225.545 148.820 1225.925 148.865 ;
        RECT 1231.045 148.820 1231.425 148.865 ;
        RECT 1225.495 148.505 1231.430 148.820 ;
        RECT 1225.545 148.485 1225.925 148.505 ;
        RECT 1231.045 148.485 1231.425 148.505 ;
        RECT 1235.045 148.485 1235.425 148.865 ;
        RECT 1239.045 148.485 1239.425 148.865 ;
        RECT 1255.980 148.395 1256.360 148.775 ;
        RECT 1259.980 148.395 1260.360 148.775 ;
        RECT 1263.980 148.730 1264.360 148.775 ;
        RECT 1269.480 148.730 1269.860 148.775 ;
        RECT 1263.930 148.415 1269.865 148.730 ;
        RECT 1263.980 148.395 1264.360 148.415 ;
        RECT 1269.480 148.395 1269.860 148.415 ;
        RECT 1273.480 148.395 1273.860 148.775 ;
        RECT 1277.480 148.395 1277.860 148.775 ;
        RECT 1283.190 148.695 1284.930 148.985 ;
        RECT 1286.980 148.645 1288.180 148.935 ;
        RECT 1289.690 148.605 1292.320 149.060 ;
        RECT 1293.900 148.710 1294.280 149.090 ;
        RECT 1198.900 148.025 1212.725 148.325 ;
        RECT 1214.400 147.860 1230.410 148.235 ;
        RECT 1248.070 147.770 1268.845 148.145 ;
        RECT 1281.470 147.935 1295.085 148.235 ;
        RECT 1198.905 147.280 1217.325 147.580 ;
        RECT 1218.770 147.270 1246.080 147.610 ;
        RECT 1257.205 147.180 1279.760 147.520 ;
        RECT 1280.870 147.190 1295.515 147.490 ;
        RECT 1198.385 146.565 1205.645 146.865 ;
        RECT 1018.060 146.140 1036.730 146.150 ;
        RECT 1018.060 146.060 1048.080 146.140 ;
        RECT 1018.060 146.050 1075.165 146.060 ;
        RECT 1018.060 145.830 1084.170 146.050 ;
        RECT 1183.440 145.945 1187.565 146.215 ;
        RECT 1198.940 146.030 1203.025 146.300 ;
        RECT 1209.345 146.265 1213.095 146.540 ;
        RECT 1214.400 146.505 1240.630 146.895 ;
        RECT 1247.100 146.415 1279.065 146.805 ;
        RECT 1291.875 146.175 1295.005 146.450 ;
        RECT 1295.750 146.415 1296.130 153.575 ;
        RECT 1296.990 151.115 1303.730 151.415 ;
        RECT 1297.580 149.320 1301.035 149.760 ;
        RECT 1304.040 149.160 1304.420 149.540 ;
        RECT 1302.440 148.645 1303.640 148.935 ;
        RECT 1309.360 148.710 1309.740 149.090 ;
        RECT 1296.395 147.935 1312.315 148.235 ;
        RECT 1296.930 147.190 1313.875 147.490 ;
        RECT 1214.400 146.140 1233.070 146.150 ;
        RECT 1214.400 146.060 1244.420 146.140 ;
        RECT 1214.400 146.050 1271.505 146.060 ;
        RECT 1214.400 145.830 1280.510 146.050 ;
        RECT 458.550 145.705 495.115 145.795 ;
        RECT 654.925 145.740 691.490 145.830 ;
        RECT 851.265 145.740 887.830 145.830 ;
        RECT 1047.605 145.740 1084.170 145.830 ;
        RECT 1243.945 145.740 1280.510 145.830 ;
        RECT 6.515 145.385 10.645 145.685 ;
        RECT -59.685 144.585 -56.120 144.595 ;
        RECT -59.685 144.260 -55.325 144.585 ;
        RECT -9.360 144.340 -3.445 144.675 ;
        RECT -6.090 144.320 -3.445 144.340 ;
        RECT -56.280 144.250 -55.325 144.260 ;
        RECT -79.090 143.620 -75.790 144.000 ;
        RECT -75.090 143.620 -71.790 144.000 ;
        RECT -65.590 143.620 -62.290 144.000 ;
        RECT -61.590 143.620 -58.290 144.000 ;
        RECT -28.765 143.700 -25.465 144.080 ;
        RECT -24.765 143.700 -21.465 144.080 ;
        RECT -15.265 143.700 -11.965 144.080 ;
        RECT -11.265 143.700 -7.965 144.080 ;
        RECT -79.090 141.620 -77.805 142.000 ;
        RECT -59.775 141.620 -58.290 142.000 ;
        RECT -28.765 141.700 -27.480 142.080 ;
        RECT -9.450 141.700 -7.965 142.080 ;
        RECT -77.585 140.940 -76.065 141.300 ;
        RECT -27.260 141.020 -25.740 141.380 ;
        RECT 4.140 139.555 4.520 145.385 ;
        RECT 13.020 145.335 17.520 145.645 ;
        RECT 21.975 145.385 26.105 145.685 ;
        RECT 8.980 144.785 15.370 145.075 ;
        RECT 8.395 144.205 19.050 144.540 ;
        RECT 7.745 143.620 10.665 143.920 ;
        RECT 14.210 143.605 17.580 143.905 ;
        RECT 5.960 142.870 6.340 143.250 ;
        RECT 8.365 142.885 10.145 143.175 ;
        RECT 11.620 142.975 12.810 143.260 ;
        RECT 15.740 142.855 17.050 143.175 ;
        RECT 7.095 142.270 7.475 142.650 ;
        RECT 10.840 142.310 11.220 142.690 ;
        RECT 13.550 142.300 13.930 142.680 ;
        RECT 14.960 142.145 18.140 142.465 ;
        RECT 4.890 139.555 8.985 139.560 ;
        RECT 19.600 139.555 19.980 145.385 ;
        RECT 28.480 145.335 32.980 145.645 ;
        RECT 119.965 145.295 124.095 145.595 ;
        RECT 35.710 145.085 71.620 145.175 ;
        RECT 24.440 144.785 30.830 145.075 ;
        RECT 35.710 144.905 102.750 145.085 ;
        RECT 71.005 144.815 102.750 144.905 ;
        RECT 106.970 144.695 113.360 144.985 ;
        RECT 23.855 144.205 34.360 144.540 ;
        RECT 59.330 144.340 69.880 144.675 ;
        RECT 106.385 144.115 116.865 144.450 ;
        RECT 23.205 143.620 26.125 143.920 ;
        RECT 29.670 143.605 33.040 143.905 ;
        RECT 37.920 143.700 39.225 144.080 ;
        RECT 39.925 143.700 43.225 144.080 ;
        RECT 43.925 143.700 47.225 144.080 ;
        RECT 47.925 143.700 49.285 144.080 ;
        RECT 51.260 143.700 52.725 144.080 ;
        RECT 53.425 143.700 56.725 144.080 ;
        RECT 57.425 143.700 60.725 144.080 ;
        RECT 61.425 143.700 62.605 144.080 ;
        RECT 76.355 143.610 77.660 143.990 ;
        RECT 82.360 143.610 85.660 143.990 ;
        RECT 86.360 143.610 87.720 143.990 ;
        RECT 89.695 143.610 91.160 143.990 ;
        RECT 91.860 143.610 95.160 143.990 ;
        RECT 99.860 143.610 101.040 143.990 ;
        RECT 39.385 143.355 39.765 143.390 ;
        RECT 21.420 142.870 21.800 143.250 ;
        RECT 23.825 142.885 25.605 143.175 ;
        RECT 27.080 142.975 28.270 143.260 ;
        RECT 31.200 142.855 32.510 143.175 ;
        RECT 39.120 143.045 42.130 143.355 ;
        RECT 39.385 143.010 39.765 143.045 ;
        RECT 43.385 143.010 44.475 143.390 ;
        RECT 47.385 143.385 47.765 143.390 ;
        RECT 44.905 143.020 47.770 143.385 ;
        RECT 52.885 143.365 53.265 143.390 ;
        RECT 52.870 143.045 55.015 143.365 ;
        RECT 47.385 143.010 47.765 143.020 ;
        RECT 52.885 143.010 53.265 143.045 ;
        RECT 55.930 143.010 57.265 143.390 ;
        RECT 60.885 143.370 61.265 143.390 ;
        RECT 58.420 143.050 61.330 143.370 ;
        RECT 77.820 143.265 78.200 143.300 ;
        RECT 60.885 143.010 61.265 143.050 ;
        RECT 77.555 142.955 80.565 143.265 ;
        RECT 77.820 142.920 78.200 142.955 ;
        RECT 81.820 142.920 82.910 143.300 ;
        RECT 85.820 143.295 86.200 143.300 ;
        RECT 83.340 142.930 86.205 143.295 ;
        RECT 91.320 143.275 91.700 143.300 ;
        RECT 91.305 142.955 93.450 143.275 ;
        RECT 85.820 142.920 86.200 142.930 ;
        RECT 91.320 142.920 91.700 142.955 ;
        RECT 94.365 142.920 95.700 143.300 ;
        RECT 99.320 143.280 99.700 143.300 ;
        RECT 96.855 142.960 99.765 143.280 ;
        RECT 99.320 142.920 99.700 142.960 ;
        RECT 103.950 142.780 104.330 143.160 ;
        RECT 106.355 142.795 108.135 143.085 ;
        RECT 109.610 142.885 110.800 143.170 ;
        RECT 113.730 142.765 115.040 143.085 ;
        RECT 22.555 142.270 22.935 142.650 ;
        RECT 26.300 142.310 26.680 142.690 ;
        RECT 29.010 142.300 29.390 142.680 ;
        RECT 30.420 142.145 33.600 142.465 ;
        RECT 105.085 142.180 105.465 142.560 ;
        RECT 108.830 142.220 109.210 142.600 ;
        RECT 111.540 142.210 111.920 142.590 ;
        RECT 37.735 141.700 39.225 142.080 ;
        RECT 39.925 141.700 41.210 142.080 ;
        RECT 59.240 141.700 60.725 142.080 ;
        RECT 61.425 141.700 62.500 142.080 ;
        RECT 112.950 142.055 116.130 142.375 ;
        RECT 76.170 141.610 77.660 141.990 ;
        RECT 99.860 141.610 100.935 141.990 ;
        RECT 39.385 141.010 40.475 141.390 ;
        RECT 41.430 141.020 42.950 141.380 ;
        RECT 43.870 141.015 56.720 141.350 ;
        RECT 60.885 141.345 61.265 141.390 ;
        RECT 60.150 141.045 61.460 141.345 ;
        RECT 60.885 141.010 61.265 141.045 ;
        RECT 77.820 140.920 78.910 141.300 ;
        RECT 79.865 140.930 81.385 141.290 ;
        RECT 82.305 140.925 95.155 141.260 ;
        RECT 99.320 141.255 99.700 141.300 ;
        RECT 98.585 140.955 99.895 141.255 ;
        RECT 99.320 140.920 99.700 140.955 ;
        RECT 36.240 140.425 69.320 140.500 ;
        RECT 36.240 140.150 101.330 140.425 ;
        RECT 68.380 140.060 101.330 140.150 ;
        RECT 103.125 140.050 107.385 140.405 ;
        RECT 20.350 139.555 24.445 139.560 ;
        RECT -82.775 138.575 -56.120 139.475 ;
        RECT -32.450 138.655 -5.795 139.555 ;
        RECT 3.770 139.550 8.985 139.555 ;
        RECT 19.230 139.550 24.445 139.555 ;
        RECT 34.690 139.550 74.940 139.555 ;
        RECT 3.770 139.465 74.940 139.550 ;
        RECT 101.330 139.465 106.975 139.470 ;
        RECT 117.590 139.465 117.970 145.295 ;
        RECT 126.470 145.245 130.970 145.555 ;
        RECT 202.880 145.385 207.010 145.685 ;
        RECT 122.430 144.695 128.820 144.985 ;
        RECT 121.845 144.115 137.865 144.450 ;
        RECT 186.810 144.350 192.725 144.685 ;
        RECT 190.080 144.330 192.725 144.350 ;
        RECT 121.195 143.530 124.115 143.830 ;
        RECT 127.660 143.515 131.030 143.815 ;
        RECT 167.405 143.710 170.705 144.090 ;
        RECT 171.405 143.710 174.705 144.090 ;
        RECT 180.905 143.710 184.205 144.090 ;
        RECT 184.905 143.710 188.205 144.090 ;
        RECT 119.410 142.780 119.790 143.160 ;
        RECT 121.815 142.795 123.595 143.085 ;
        RECT 125.070 142.885 126.260 143.170 ;
        RECT 129.190 142.765 130.500 143.085 ;
        RECT 120.545 142.180 120.925 142.560 ;
        RECT 124.290 142.220 124.670 142.600 ;
        RECT 127.000 142.210 127.380 142.590 ;
        RECT 128.410 142.055 131.590 142.375 ;
        RECT 167.405 141.710 168.690 142.090 ;
        RECT 186.720 141.710 188.205 142.090 ;
        RECT 118.690 140.970 122.840 141.240 ;
        RECT 168.910 141.030 170.430 141.390 ;
        RECT 118.340 139.465 122.435 139.470 ;
        RECT 3.770 139.460 106.975 139.465 ;
        RECT 117.220 139.460 122.435 139.465 ;
        RECT 3.770 138.655 132.250 139.460 ;
        RECT 163.720 138.665 190.375 139.565 ;
        RECT 200.505 139.555 200.885 145.385 ;
        RECT 209.385 145.335 213.885 145.645 ;
        RECT 218.340 145.385 222.470 145.685 ;
        RECT 205.345 144.785 211.735 145.075 ;
        RECT 204.760 144.205 215.415 144.540 ;
        RECT 204.110 143.620 207.030 143.920 ;
        RECT 210.575 143.605 213.945 143.905 ;
        RECT 202.325 142.870 202.705 143.250 ;
        RECT 204.730 142.885 206.510 143.175 ;
        RECT 207.985 142.975 209.175 143.260 ;
        RECT 212.105 142.855 213.415 143.175 ;
        RECT 203.460 142.270 203.840 142.650 ;
        RECT 207.205 142.310 207.585 142.690 ;
        RECT 209.915 142.300 210.295 142.680 ;
        RECT 211.325 142.145 214.505 142.465 ;
        RECT 201.255 139.555 205.350 139.560 ;
        RECT 215.965 139.555 216.345 145.385 ;
        RECT 224.845 145.335 229.345 145.645 ;
        RECT 316.330 145.295 320.460 145.595 ;
        RECT 232.075 145.085 267.985 145.175 ;
        RECT 220.805 144.785 227.195 145.075 ;
        RECT 232.075 144.905 299.115 145.085 ;
        RECT 267.370 144.815 299.115 144.905 ;
        RECT 303.335 144.695 309.725 144.985 ;
        RECT 220.220 144.205 230.725 144.540 ;
        RECT 255.695 144.340 266.245 144.675 ;
        RECT 302.750 144.115 313.230 144.450 ;
        RECT 219.570 143.620 222.490 143.920 ;
        RECT 226.035 143.605 229.405 143.905 ;
        RECT 234.285 143.700 235.590 144.080 ;
        RECT 236.290 143.700 239.590 144.080 ;
        RECT 240.290 143.700 243.590 144.080 ;
        RECT 244.290 143.700 245.650 144.080 ;
        RECT 247.625 143.700 249.090 144.080 ;
        RECT 249.790 143.700 253.090 144.080 ;
        RECT 253.790 143.700 257.090 144.080 ;
        RECT 257.790 143.700 258.970 144.080 ;
        RECT 272.720 143.610 274.025 143.990 ;
        RECT 278.725 143.610 282.025 143.990 ;
        RECT 282.725 143.610 284.085 143.990 ;
        RECT 286.060 143.610 287.525 143.990 ;
        RECT 288.225 143.610 291.525 143.990 ;
        RECT 296.225 143.610 297.405 143.990 ;
        RECT 235.750 143.355 236.130 143.390 ;
        RECT 217.785 142.870 218.165 143.250 ;
        RECT 220.190 142.885 221.970 143.175 ;
        RECT 223.445 142.975 224.635 143.260 ;
        RECT 227.565 142.855 228.875 143.175 ;
        RECT 235.485 143.045 238.495 143.355 ;
        RECT 235.750 143.010 236.130 143.045 ;
        RECT 239.750 143.010 240.840 143.390 ;
        RECT 243.750 143.385 244.130 143.390 ;
        RECT 241.270 143.020 244.135 143.385 ;
        RECT 249.250 143.365 249.630 143.390 ;
        RECT 249.235 143.045 251.380 143.365 ;
        RECT 243.750 143.010 244.130 143.020 ;
        RECT 249.250 143.010 249.630 143.045 ;
        RECT 252.295 143.010 253.630 143.390 ;
        RECT 257.250 143.370 257.630 143.390 ;
        RECT 254.785 143.050 257.695 143.370 ;
        RECT 274.185 143.265 274.565 143.300 ;
        RECT 257.250 143.010 257.630 143.050 ;
        RECT 273.920 142.955 276.930 143.265 ;
        RECT 274.185 142.920 274.565 142.955 ;
        RECT 278.185 142.920 279.275 143.300 ;
        RECT 282.185 143.295 282.565 143.300 ;
        RECT 279.705 142.930 282.570 143.295 ;
        RECT 287.685 143.275 288.065 143.300 ;
        RECT 287.670 142.955 289.815 143.275 ;
        RECT 282.185 142.920 282.565 142.930 ;
        RECT 287.685 142.920 288.065 142.955 ;
        RECT 290.730 142.920 292.065 143.300 ;
        RECT 295.685 143.280 296.065 143.300 ;
        RECT 293.220 142.960 296.130 143.280 ;
        RECT 295.685 142.920 296.065 142.960 ;
        RECT 300.315 142.780 300.695 143.160 ;
        RECT 302.720 142.795 304.500 143.085 ;
        RECT 305.975 142.885 307.165 143.170 ;
        RECT 310.095 142.765 311.405 143.085 ;
        RECT 218.920 142.270 219.300 142.650 ;
        RECT 222.665 142.310 223.045 142.690 ;
        RECT 225.375 142.300 225.755 142.680 ;
        RECT 226.785 142.145 229.965 142.465 ;
        RECT 301.450 142.180 301.830 142.560 ;
        RECT 305.195 142.220 305.575 142.600 ;
        RECT 307.905 142.210 308.285 142.590 ;
        RECT 234.100 141.700 235.590 142.080 ;
        RECT 236.290 141.700 237.575 142.080 ;
        RECT 255.605 141.700 257.090 142.080 ;
        RECT 257.790 141.700 258.865 142.080 ;
        RECT 309.315 142.055 312.495 142.375 ;
        RECT 272.535 141.610 274.025 141.990 ;
        RECT 296.225 141.610 297.300 141.990 ;
        RECT 235.750 141.010 236.840 141.390 ;
        RECT 237.795 141.020 239.315 141.380 ;
        RECT 240.235 141.015 253.085 141.350 ;
        RECT 257.250 141.345 257.630 141.390 ;
        RECT 256.515 141.045 257.825 141.345 ;
        RECT 257.250 141.010 257.630 141.045 ;
        RECT 274.185 140.920 275.275 141.300 ;
        RECT 276.230 140.930 277.750 141.290 ;
        RECT 278.670 140.925 291.520 141.260 ;
        RECT 295.685 141.255 296.065 141.300 ;
        RECT 294.950 140.955 296.260 141.255 ;
        RECT 295.685 140.920 296.065 140.955 ;
        RECT 232.605 140.425 265.685 140.500 ;
        RECT 232.605 140.150 297.695 140.425 ;
        RECT 264.745 140.060 297.695 140.150 ;
        RECT 299.490 140.050 303.750 140.405 ;
        RECT 216.715 139.555 220.810 139.560 ;
        RECT 200.135 139.550 205.350 139.555 ;
        RECT 215.595 139.550 220.810 139.555 ;
        RECT 231.055 139.550 271.305 139.555 ;
        RECT 200.135 139.465 271.305 139.550 ;
        RECT 297.695 139.465 303.340 139.470 ;
        RECT 313.955 139.465 314.335 145.295 ;
        RECT 322.835 145.245 327.335 145.555 ;
        RECT 399.280 145.335 403.410 145.635 ;
        RECT 318.795 144.695 325.185 144.985 ;
        RECT 318.210 144.115 334.230 144.450 ;
        RECT 383.200 144.310 389.115 144.645 ;
        RECT 386.470 144.290 389.115 144.310 ;
        RECT 317.560 143.530 320.480 143.830 ;
        RECT 324.025 143.515 327.395 143.815 ;
        RECT 363.795 143.670 367.095 144.050 ;
        RECT 367.795 143.670 371.095 144.050 ;
        RECT 377.295 143.670 380.595 144.050 ;
        RECT 381.295 143.670 384.595 144.050 ;
        RECT 315.775 142.780 316.155 143.160 ;
        RECT 318.180 142.795 319.960 143.085 ;
        RECT 321.435 142.885 322.625 143.170 ;
        RECT 325.555 142.765 326.865 143.085 ;
        RECT 316.910 142.180 317.290 142.560 ;
        RECT 320.655 142.220 321.035 142.600 ;
        RECT 323.365 142.210 323.745 142.590 ;
        RECT 324.775 142.055 327.955 142.375 ;
        RECT 363.795 141.670 365.080 142.050 ;
        RECT 383.110 141.670 384.595 142.050 ;
        RECT 315.055 140.970 319.205 141.240 ;
        RECT 365.300 140.990 366.820 141.350 ;
        RECT 314.705 139.465 318.800 139.470 ;
        RECT 200.135 139.460 303.340 139.465 ;
        RECT 313.585 139.460 318.800 139.465 ;
        RECT 200.135 138.655 328.615 139.460 ;
        RECT 74.675 138.565 132.250 138.655 ;
        RECT 271.040 138.565 328.615 138.655 ;
        RECT 360.110 138.625 386.765 139.525 ;
        RECT 396.905 139.505 397.285 145.335 ;
        RECT 405.785 145.285 410.285 145.595 ;
        RECT 414.740 145.335 418.870 145.635 ;
        RECT 401.745 144.735 408.135 145.025 ;
        RECT 401.160 144.155 411.815 144.490 ;
        RECT 400.510 143.570 403.430 143.870 ;
        RECT 406.975 143.555 410.345 143.855 ;
        RECT 398.725 142.820 399.105 143.200 ;
        RECT 401.130 142.835 402.910 143.125 ;
        RECT 404.385 142.925 405.575 143.210 ;
        RECT 408.505 142.805 409.815 143.125 ;
        RECT 399.860 142.220 400.240 142.600 ;
        RECT 403.605 142.260 403.985 142.640 ;
        RECT 406.315 142.250 406.695 142.630 ;
        RECT 407.725 142.095 410.905 142.415 ;
        RECT 397.655 139.505 401.750 139.510 ;
        RECT 412.365 139.505 412.745 145.335 ;
        RECT 421.245 145.285 425.745 145.595 ;
        RECT 512.730 145.245 516.860 145.545 ;
        RECT 428.475 145.035 464.385 145.125 ;
        RECT 417.205 144.735 423.595 145.025 ;
        RECT 428.475 144.855 495.515 145.035 ;
        RECT 463.770 144.765 495.515 144.855 ;
        RECT 499.735 144.645 506.125 144.935 ;
        RECT 416.620 144.155 427.125 144.490 ;
        RECT 452.095 144.290 462.645 144.625 ;
        RECT 499.150 144.065 509.630 144.400 ;
        RECT 415.970 143.570 418.890 143.870 ;
        RECT 422.435 143.555 425.805 143.855 ;
        RECT 430.685 143.650 431.990 144.030 ;
        RECT 432.690 143.650 435.990 144.030 ;
        RECT 436.690 143.650 439.990 144.030 ;
        RECT 440.690 143.650 442.050 144.030 ;
        RECT 444.025 143.650 445.490 144.030 ;
        RECT 446.190 143.650 449.490 144.030 ;
        RECT 450.190 143.650 453.490 144.030 ;
        RECT 454.190 143.650 455.370 144.030 ;
        RECT 469.120 143.560 470.425 143.940 ;
        RECT 475.125 143.560 478.425 143.940 ;
        RECT 479.125 143.560 480.485 143.940 ;
        RECT 482.460 143.560 483.925 143.940 ;
        RECT 484.625 143.560 487.925 143.940 ;
        RECT 492.625 143.560 493.805 143.940 ;
        RECT 432.150 143.305 432.530 143.340 ;
        RECT 414.185 142.820 414.565 143.200 ;
        RECT 416.590 142.835 418.370 143.125 ;
        RECT 419.845 142.925 421.035 143.210 ;
        RECT 423.965 142.805 425.275 143.125 ;
        RECT 431.885 142.995 434.895 143.305 ;
        RECT 432.150 142.960 432.530 142.995 ;
        RECT 436.150 142.960 437.240 143.340 ;
        RECT 440.150 143.335 440.530 143.340 ;
        RECT 437.670 142.970 440.535 143.335 ;
        RECT 445.650 143.315 446.030 143.340 ;
        RECT 445.635 142.995 447.780 143.315 ;
        RECT 440.150 142.960 440.530 142.970 ;
        RECT 445.650 142.960 446.030 142.995 ;
        RECT 448.695 142.960 450.030 143.340 ;
        RECT 453.650 143.320 454.030 143.340 ;
        RECT 451.185 143.000 454.095 143.320 ;
        RECT 470.585 143.215 470.965 143.250 ;
        RECT 453.650 142.960 454.030 143.000 ;
        RECT 470.320 142.905 473.330 143.215 ;
        RECT 470.585 142.870 470.965 142.905 ;
        RECT 474.585 142.870 475.675 143.250 ;
        RECT 478.585 143.245 478.965 143.250 ;
        RECT 476.105 142.880 478.970 143.245 ;
        RECT 484.085 143.225 484.465 143.250 ;
        RECT 484.070 142.905 486.215 143.225 ;
        RECT 478.585 142.870 478.965 142.880 ;
        RECT 484.085 142.870 484.465 142.905 ;
        RECT 487.130 142.870 488.465 143.250 ;
        RECT 492.085 143.230 492.465 143.250 ;
        RECT 489.620 142.910 492.530 143.230 ;
        RECT 492.085 142.870 492.465 142.910 ;
        RECT 496.715 142.730 497.095 143.110 ;
        RECT 499.120 142.745 500.900 143.035 ;
        RECT 502.375 142.835 503.565 143.120 ;
        RECT 506.495 142.715 507.805 143.035 ;
        RECT 415.320 142.220 415.700 142.600 ;
        RECT 419.065 142.260 419.445 142.640 ;
        RECT 421.775 142.250 422.155 142.630 ;
        RECT 423.185 142.095 426.365 142.415 ;
        RECT 497.850 142.130 498.230 142.510 ;
        RECT 501.595 142.170 501.975 142.550 ;
        RECT 504.305 142.160 504.685 142.540 ;
        RECT 430.500 141.650 431.990 142.030 ;
        RECT 432.690 141.650 433.975 142.030 ;
        RECT 452.005 141.650 453.490 142.030 ;
        RECT 454.190 141.650 455.265 142.030 ;
        RECT 505.715 142.005 508.895 142.325 ;
        RECT 468.935 141.560 470.425 141.940 ;
        RECT 492.625 141.560 493.700 141.940 ;
        RECT 432.150 140.960 433.240 141.340 ;
        RECT 434.195 140.970 435.715 141.330 ;
        RECT 436.635 140.965 449.485 141.300 ;
        RECT 453.650 141.295 454.030 141.340 ;
        RECT 452.915 140.995 454.225 141.295 ;
        RECT 453.650 140.960 454.030 140.995 ;
        RECT 470.585 140.870 471.675 141.250 ;
        RECT 472.630 140.880 474.150 141.240 ;
        RECT 475.070 140.875 487.920 141.210 ;
        RECT 492.085 141.205 492.465 141.250 ;
        RECT 491.350 140.905 492.660 141.205 ;
        RECT 492.085 140.870 492.465 140.905 ;
        RECT 429.005 140.375 462.085 140.450 ;
        RECT 429.005 140.100 494.095 140.375 ;
        RECT 461.145 140.010 494.095 140.100 ;
        RECT 495.890 140.000 500.150 140.355 ;
        RECT 413.115 139.505 417.210 139.510 ;
        RECT 396.535 139.500 401.750 139.505 ;
        RECT 411.995 139.500 417.210 139.505 ;
        RECT 427.455 139.500 467.705 139.505 ;
        RECT 396.535 139.415 467.705 139.500 ;
        RECT 494.095 139.415 499.740 139.420 ;
        RECT 510.355 139.415 510.735 145.245 ;
        RECT 519.235 145.195 523.735 145.505 ;
        RECT 595.655 145.370 599.785 145.670 ;
        RECT 515.195 144.645 521.585 144.935 ;
        RECT 514.610 144.065 530.630 144.400 ;
        RECT 579.520 144.355 585.435 144.690 ;
        RECT 582.790 144.335 585.435 144.355 ;
        RECT 513.960 143.480 516.880 143.780 ;
        RECT 520.425 143.465 523.795 143.765 ;
        RECT 560.115 143.715 563.415 144.095 ;
        RECT 564.115 143.715 567.415 144.095 ;
        RECT 573.615 143.715 576.915 144.095 ;
        RECT 577.615 143.715 580.915 144.095 ;
        RECT 512.175 142.730 512.555 143.110 ;
        RECT 514.580 142.745 516.360 143.035 ;
        RECT 517.835 142.835 519.025 143.120 ;
        RECT 521.955 142.715 523.265 143.035 ;
        RECT 513.310 142.130 513.690 142.510 ;
        RECT 517.055 142.170 517.435 142.550 ;
        RECT 519.765 142.160 520.145 142.540 ;
        RECT 521.175 142.005 524.355 142.325 ;
        RECT 560.115 141.715 561.400 142.095 ;
        RECT 579.430 141.715 580.915 142.095 ;
        RECT 511.455 140.920 515.605 141.190 ;
        RECT 561.620 141.035 563.140 141.395 ;
        RECT 511.105 139.415 515.200 139.420 ;
        RECT 396.535 139.410 499.740 139.415 ;
        RECT 509.985 139.410 515.200 139.415 ;
        RECT 396.535 138.605 525.015 139.410 ;
        RECT 556.430 138.670 583.085 139.570 ;
        RECT 593.280 139.540 593.660 145.370 ;
        RECT 602.160 145.320 606.660 145.630 ;
        RECT 611.115 145.370 615.245 145.670 ;
        RECT 598.120 144.770 604.510 145.060 ;
        RECT 597.535 144.190 608.190 144.525 ;
        RECT 596.885 143.605 599.805 143.905 ;
        RECT 603.350 143.590 606.720 143.890 ;
        RECT 595.100 142.855 595.480 143.235 ;
        RECT 597.505 142.870 599.285 143.160 ;
        RECT 600.760 142.960 601.950 143.245 ;
        RECT 604.880 142.840 606.190 143.160 ;
        RECT 596.235 142.255 596.615 142.635 ;
        RECT 599.980 142.295 600.360 142.675 ;
        RECT 602.690 142.285 603.070 142.665 ;
        RECT 604.100 142.130 607.280 142.450 ;
        RECT 594.030 139.540 598.125 139.545 ;
        RECT 608.740 139.540 609.120 145.370 ;
        RECT 617.620 145.320 622.120 145.630 ;
        RECT 709.105 145.280 713.235 145.580 ;
        RECT 624.850 145.070 660.760 145.160 ;
        RECT 613.580 144.770 619.970 145.060 ;
        RECT 624.850 144.890 691.890 145.070 ;
        RECT 660.145 144.800 691.890 144.890 ;
        RECT 696.110 144.680 702.500 144.970 ;
        RECT 612.995 144.190 623.500 144.525 ;
        RECT 648.470 144.325 659.020 144.660 ;
        RECT 695.525 144.100 706.005 144.435 ;
        RECT 612.345 143.605 615.265 143.905 ;
        RECT 618.810 143.590 622.180 143.890 ;
        RECT 627.060 143.685 628.365 144.065 ;
        RECT 629.065 143.685 632.365 144.065 ;
        RECT 633.065 143.685 636.365 144.065 ;
        RECT 637.065 143.685 638.425 144.065 ;
        RECT 640.400 143.685 641.865 144.065 ;
        RECT 642.565 143.685 645.865 144.065 ;
        RECT 646.565 143.685 649.865 144.065 ;
        RECT 650.565 143.685 651.745 144.065 ;
        RECT 665.495 143.595 666.800 143.975 ;
        RECT 671.500 143.595 674.800 143.975 ;
        RECT 675.500 143.595 676.860 143.975 ;
        RECT 678.835 143.595 680.300 143.975 ;
        RECT 681.000 143.595 684.300 143.975 ;
        RECT 689.000 143.595 690.180 143.975 ;
        RECT 628.525 143.340 628.905 143.375 ;
        RECT 610.560 142.855 610.940 143.235 ;
        RECT 612.965 142.870 614.745 143.160 ;
        RECT 616.220 142.960 617.410 143.245 ;
        RECT 620.340 142.840 621.650 143.160 ;
        RECT 628.260 143.030 631.270 143.340 ;
        RECT 628.525 142.995 628.905 143.030 ;
        RECT 632.525 142.995 633.615 143.375 ;
        RECT 636.525 143.370 636.905 143.375 ;
        RECT 634.045 143.005 636.910 143.370 ;
        RECT 642.025 143.350 642.405 143.375 ;
        RECT 642.010 143.030 644.155 143.350 ;
        RECT 636.525 142.995 636.905 143.005 ;
        RECT 642.025 142.995 642.405 143.030 ;
        RECT 645.070 142.995 646.405 143.375 ;
        RECT 650.025 143.355 650.405 143.375 ;
        RECT 647.560 143.035 650.470 143.355 ;
        RECT 666.960 143.250 667.340 143.285 ;
        RECT 650.025 142.995 650.405 143.035 ;
        RECT 666.695 142.940 669.705 143.250 ;
        RECT 666.960 142.905 667.340 142.940 ;
        RECT 670.960 142.905 672.050 143.285 ;
        RECT 674.960 143.280 675.340 143.285 ;
        RECT 672.480 142.915 675.345 143.280 ;
        RECT 680.460 143.260 680.840 143.285 ;
        RECT 680.445 142.940 682.590 143.260 ;
        RECT 674.960 142.905 675.340 142.915 ;
        RECT 680.460 142.905 680.840 142.940 ;
        RECT 683.505 142.905 684.840 143.285 ;
        RECT 688.460 143.265 688.840 143.285 ;
        RECT 685.995 142.945 688.905 143.265 ;
        RECT 688.460 142.905 688.840 142.945 ;
        RECT 693.090 142.765 693.470 143.145 ;
        RECT 695.495 142.780 697.275 143.070 ;
        RECT 698.750 142.870 699.940 143.155 ;
        RECT 702.870 142.750 704.180 143.070 ;
        RECT 611.695 142.255 612.075 142.635 ;
        RECT 615.440 142.295 615.820 142.675 ;
        RECT 618.150 142.285 618.530 142.665 ;
        RECT 619.560 142.130 622.740 142.450 ;
        RECT 694.225 142.165 694.605 142.545 ;
        RECT 697.970 142.205 698.350 142.585 ;
        RECT 700.680 142.195 701.060 142.575 ;
        RECT 626.875 141.685 628.365 142.065 ;
        RECT 629.065 141.685 630.350 142.065 ;
        RECT 648.380 141.685 649.865 142.065 ;
        RECT 650.565 141.685 651.640 142.065 ;
        RECT 702.090 142.040 705.270 142.360 ;
        RECT 665.310 141.595 666.800 141.975 ;
        RECT 689.000 141.595 690.075 141.975 ;
        RECT 628.525 140.995 629.615 141.375 ;
        RECT 630.570 141.005 632.090 141.365 ;
        RECT 633.010 141.000 645.860 141.335 ;
        RECT 650.025 141.330 650.405 141.375 ;
        RECT 649.290 141.030 650.600 141.330 ;
        RECT 650.025 140.995 650.405 141.030 ;
        RECT 666.960 140.905 668.050 141.285 ;
        RECT 669.005 140.915 670.525 141.275 ;
        RECT 671.445 140.910 684.295 141.245 ;
        RECT 688.460 141.240 688.840 141.285 ;
        RECT 687.725 140.940 689.035 141.240 ;
        RECT 688.460 140.905 688.840 140.940 ;
        RECT 625.380 140.410 658.460 140.485 ;
        RECT 625.380 140.135 690.470 140.410 ;
        RECT 657.520 140.045 690.470 140.135 ;
        RECT 692.265 140.035 696.525 140.390 ;
        RECT 609.490 139.540 613.585 139.545 ;
        RECT 592.910 139.535 598.125 139.540 ;
        RECT 608.370 139.535 613.585 139.540 ;
        RECT 623.830 139.535 664.080 139.540 ;
        RECT 592.910 139.450 664.080 139.535 ;
        RECT 690.470 139.450 696.115 139.455 ;
        RECT 706.730 139.450 707.110 145.280 ;
        RECT 715.610 145.230 720.110 145.540 ;
        RECT 791.995 145.370 796.125 145.670 ;
        RECT 711.570 144.680 717.960 144.970 ;
        RECT 710.985 144.100 727.005 144.435 ;
        RECT 775.885 144.360 781.800 144.695 ;
        RECT 779.155 144.340 781.800 144.360 ;
        RECT 710.335 143.515 713.255 143.815 ;
        RECT 716.800 143.500 720.170 143.800 ;
        RECT 756.480 143.720 759.780 144.100 ;
        RECT 760.480 143.720 763.780 144.100 ;
        RECT 769.980 143.720 773.280 144.100 ;
        RECT 773.980 143.720 777.280 144.100 ;
        RECT 708.550 142.765 708.930 143.145 ;
        RECT 710.955 142.780 712.735 143.070 ;
        RECT 714.210 142.870 715.400 143.155 ;
        RECT 718.330 142.750 719.640 143.070 ;
        RECT 709.685 142.165 710.065 142.545 ;
        RECT 713.430 142.205 713.810 142.585 ;
        RECT 716.140 142.195 716.520 142.575 ;
        RECT 717.550 142.040 720.730 142.360 ;
        RECT 756.480 141.720 757.765 142.100 ;
        RECT 775.795 141.720 777.280 142.100 ;
        RECT 707.830 140.955 711.980 141.225 ;
        RECT 757.985 141.040 759.505 141.400 ;
        RECT 707.480 139.450 711.575 139.455 ;
        RECT 592.910 139.445 696.115 139.450 ;
        RECT 706.360 139.445 711.575 139.450 ;
        RECT 592.910 138.640 721.390 139.445 ;
        RECT 752.795 138.675 779.450 139.575 ;
        RECT 789.620 139.540 790.000 145.370 ;
        RECT 798.500 145.320 803.000 145.630 ;
        RECT 807.455 145.370 811.585 145.670 ;
        RECT 794.460 144.770 800.850 145.060 ;
        RECT 793.875 144.190 804.530 144.525 ;
        RECT 793.225 143.605 796.145 143.905 ;
        RECT 799.690 143.590 803.060 143.890 ;
        RECT 791.440 142.855 791.820 143.235 ;
        RECT 793.845 142.870 795.625 143.160 ;
        RECT 797.100 142.960 798.290 143.245 ;
        RECT 801.220 142.840 802.530 143.160 ;
        RECT 792.575 142.255 792.955 142.635 ;
        RECT 796.320 142.295 796.700 142.675 ;
        RECT 799.030 142.285 799.410 142.665 ;
        RECT 800.440 142.130 803.620 142.450 ;
        RECT 790.370 139.540 794.465 139.545 ;
        RECT 805.080 139.540 805.460 145.370 ;
        RECT 813.960 145.320 818.460 145.630 ;
        RECT 905.445 145.280 909.575 145.580 ;
        RECT 821.190 145.070 857.100 145.160 ;
        RECT 809.920 144.770 816.310 145.060 ;
        RECT 821.190 144.890 888.230 145.070 ;
        RECT 856.485 144.800 888.230 144.890 ;
        RECT 892.450 144.680 898.840 144.970 ;
        RECT 809.335 144.190 819.840 144.525 ;
        RECT 844.810 144.325 855.360 144.660 ;
        RECT 891.865 144.100 902.345 144.435 ;
        RECT 808.685 143.605 811.605 143.905 ;
        RECT 815.150 143.590 818.520 143.890 ;
        RECT 823.400 143.685 824.705 144.065 ;
        RECT 825.405 143.685 828.705 144.065 ;
        RECT 829.405 143.685 832.705 144.065 ;
        RECT 833.405 143.685 834.765 144.065 ;
        RECT 836.740 143.685 838.205 144.065 ;
        RECT 838.905 143.685 842.205 144.065 ;
        RECT 842.905 143.685 846.205 144.065 ;
        RECT 846.905 143.685 848.085 144.065 ;
        RECT 861.835 143.595 863.140 143.975 ;
        RECT 867.840 143.595 871.140 143.975 ;
        RECT 871.840 143.595 873.200 143.975 ;
        RECT 875.175 143.595 876.640 143.975 ;
        RECT 877.340 143.595 880.640 143.975 ;
        RECT 885.340 143.595 886.520 143.975 ;
        RECT 824.865 143.340 825.245 143.375 ;
        RECT 806.900 142.855 807.280 143.235 ;
        RECT 809.305 142.870 811.085 143.160 ;
        RECT 812.560 142.960 813.750 143.245 ;
        RECT 816.680 142.840 817.990 143.160 ;
        RECT 824.600 143.030 827.610 143.340 ;
        RECT 824.865 142.995 825.245 143.030 ;
        RECT 828.865 142.995 829.955 143.375 ;
        RECT 832.865 143.370 833.245 143.375 ;
        RECT 830.385 143.005 833.250 143.370 ;
        RECT 838.365 143.350 838.745 143.375 ;
        RECT 838.350 143.030 840.495 143.350 ;
        RECT 832.865 142.995 833.245 143.005 ;
        RECT 838.365 142.995 838.745 143.030 ;
        RECT 841.410 142.995 842.745 143.375 ;
        RECT 846.365 143.355 846.745 143.375 ;
        RECT 843.900 143.035 846.810 143.355 ;
        RECT 863.300 143.250 863.680 143.285 ;
        RECT 846.365 142.995 846.745 143.035 ;
        RECT 863.035 142.940 866.045 143.250 ;
        RECT 863.300 142.905 863.680 142.940 ;
        RECT 867.300 142.905 868.390 143.285 ;
        RECT 871.300 143.280 871.680 143.285 ;
        RECT 868.820 142.915 871.685 143.280 ;
        RECT 876.800 143.260 877.180 143.285 ;
        RECT 876.785 142.940 878.930 143.260 ;
        RECT 871.300 142.905 871.680 142.915 ;
        RECT 876.800 142.905 877.180 142.940 ;
        RECT 879.845 142.905 881.180 143.285 ;
        RECT 884.800 143.265 885.180 143.285 ;
        RECT 882.335 142.945 885.245 143.265 ;
        RECT 884.800 142.905 885.180 142.945 ;
        RECT 889.430 142.765 889.810 143.145 ;
        RECT 891.835 142.780 893.615 143.070 ;
        RECT 895.090 142.870 896.280 143.155 ;
        RECT 899.210 142.750 900.520 143.070 ;
        RECT 808.035 142.255 808.415 142.635 ;
        RECT 811.780 142.295 812.160 142.675 ;
        RECT 814.490 142.285 814.870 142.665 ;
        RECT 815.900 142.130 819.080 142.450 ;
        RECT 890.565 142.165 890.945 142.545 ;
        RECT 894.310 142.205 894.690 142.585 ;
        RECT 897.020 142.195 897.400 142.575 ;
        RECT 823.215 141.685 824.705 142.065 ;
        RECT 825.405 141.685 826.690 142.065 ;
        RECT 844.720 141.685 846.205 142.065 ;
        RECT 846.905 141.685 847.980 142.065 ;
        RECT 898.430 142.040 901.610 142.360 ;
        RECT 861.650 141.595 863.140 141.975 ;
        RECT 885.340 141.595 886.415 141.975 ;
        RECT 824.865 140.995 825.955 141.375 ;
        RECT 826.910 141.005 828.430 141.365 ;
        RECT 829.350 141.000 842.200 141.335 ;
        RECT 846.365 141.330 846.745 141.375 ;
        RECT 845.630 141.030 846.940 141.330 ;
        RECT 846.365 140.995 846.745 141.030 ;
        RECT 863.300 140.905 864.390 141.285 ;
        RECT 865.345 140.915 866.865 141.275 ;
        RECT 867.785 140.910 880.635 141.245 ;
        RECT 884.800 141.240 885.180 141.285 ;
        RECT 884.065 140.940 885.375 141.240 ;
        RECT 884.800 140.905 885.180 140.940 ;
        RECT 821.720 140.410 854.800 140.485 ;
        RECT 821.720 140.135 886.810 140.410 ;
        RECT 853.860 140.045 886.810 140.135 ;
        RECT 888.605 140.035 892.865 140.390 ;
        RECT 805.830 139.540 809.925 139.545 ;
        RECT 789.250 139.535 794.465 139.540 ;
        RECT 804.710 139.535 809.925 139.540 ;
        RECT 820.170 139.535 860.420 139.540 ;
        RECT 789.250 139.450 860.420 139.535 ;
        RECT 886.810 139.450 892.455 139.455 ;
        RECT 903.070 139.450 903.450 145.280 ;
        RECT 911.950 145.230 916.450 145.540 ;
        RECT 988.335 145.370 992.465 145.670 ;
        RECT 907.910 144.680 914.300 144.970 ;
        RECT 907.325 144.100 923.345 144.435 ;
        RECT 972.270 144.345 978.185 144.680 ;
        RECT 975.540 144.325 978.185 144.345 ;
        RECT 906.675 143.515 909.595 143.815 ;
        RECT 913.140 143.500 916.510 143.800 ;
        RECT 952.865 143.705 956.165 144.085 ;
        RECT 956.865 143.705 960.165 144.085 ;
        RECT 966.365 143.705 969.665 144.085 ;
        RECT 970.365 143.705 973.665 144.085 ;
        RECT 904.890 142.765 905.270 143.145 ;
        RECT 907.295 142.780 909.075 143.070 ;
        RECT 910.550 142.870 911.740 143.155 ;
        RECT 914.670 142.750 915.980 143.070 ;
        RECT 906.025 142.165 906.405 142.545 ;
        RECT 909.770 142.205 910.150 142.585 ;
        RECT 912.480 142.195 912.860 142.575 ;
        RECT 913.890 142.040 917.070 142.360 ;
        RECT 952.865 141.705 954.150 142.085 ;
        RECT 972.180 141.705 973.665 142.085 ;
        RECT 904.170 140.955 908.320 141.225 ;
        RECT 954.370 141.025 955.890 141.385 ;
        RECT 903.820 139.450 907.915 139.455 ;
        RECT 789.250 139.445 892.455 139.450 ;
        RECT 902.700 139.445 907.915 139.450 ;
        RECT 789.250 138.640 917.730 139.445 ;
        RECT 949.180 138.660 975.835 139.560 ;
        RECT 985.960 139.540 986.340 145.370 ;
        RECT 994.840 145.320 999.340 145.630 ;
        RECT 1003.795 145.370 1007.925 145.670 ;
        RECT 990.800 144.770 997.190 145.060 ;
        RECT 990.215 144.190 1000.870 144.525 ;
        RECT 989.565 143.605 992.485 143.905 ;
        RECT 996.030 143.590 999.400 143.890 ;
        RECT 987.780 142.855 988.160 143.235 ;
        RECT 990.185 142.870 991.965 143.160 ;
        RECT 993.440 142.960 994.630 143.245 ;
        RECT 997.560 142.840 998.870 143.160 ;
        RECT 988.915 142.255 989.295 142.635 ;
        RECT 992.660 142.295 993.040 142.675 ;
        RECT 995.370 142.285 995.750 142.665 ;
        RECT 996.780 142.130 999.960 142.450 ;
        RECT 986.710 139.540 990.805 139.545 ;
        RECT 1001.420 139.540 1001.800 145.370 ;
        RECT 1010.300 145.320 1014.800 145.630 ;
        RECT 1101.785 145.280 1105.915 145.580 ;
        RECT 1017.530 145.070 1053.440 145.160 ;
        RECT 1006.260 144.770 1012.650 145.060 ;
        RECT 1017.530 144.890 1084.570 145.070 ;
        RECT 1052.825 144.800 1084.570 144.890 ;
        RECT 1088.790 144.680 1095.180 144.970 ;
        RECT 1005.675 144.190 1016.180 144.525 ;
        RECT 1041.150 144.325 1051.700 144.660 ;
        RECT 1088.205 144.100 1098.685 144.435 ;
        RECT 1005.025 143.605 1007.945 143.905 ;
        RECT 1011.490 143.590 1014.860 143.890 ;
        RECT 1019.740 143.685 1021.045 144.065 ;
        RECT 1021.745 143.685 1025.045 144.065 ;
        RECT 1025.745 143.685 1029.045 144.065 ;
        RECT 1029.745 143.685 1031.105 144.065 ;
        RECT 1033.080 143.685 1034.545 144.065 ;
        RECT 1035.245 143.685 1038.545 144.065 ;
        RECT 1039.245 143.685 1042.545 144.065 ;
        RECT 1043.245 143.685 1044.425 144.065 ;
        RECT 1058.175 143.595 1059.480 143.975 ;
        RECT 1064.180 143.595 1067.480 143.975 ;
        RECT 1068.180 143.595 1069.540 143.975 ;
        RECT 1071.515 143.595 1072.980 143.975 ;
        RECT 1073.680 143.595 1076.980 143.975 ;
        RECT 1081.680 143.595 1082.860 143.975 ;
        RECT 1021.205 143.340 1021.585 143.375 ;
        RECT 1003.240 142.855 1003.620 143.235 ;
        RECT 1005.645 142.870 1007.425 143.160 ;
        RECT 1008.900 142.960 1010.090 143.245 ;
        RECT 1013.020 142.840 1014.330 143.160 ;
        RECT 1020.940 143.030 1023.950 143.340 ;
        RECT 1021.205 142.995 1021.585 143.030 ;
        RECT 1025.205 142.995 1026.295 143.375 ;
        RECT 1029.205 143.370 1029.585 143.375 ;
        RECT 1026.725 143.005 1029.590 143.370 ;
        RECT 1034.705 143.350 1035.085 143.375 ;
        RECT 1034.690 143.030 1036.835 143.350 ;
        RECT 1029.205 142.995 1029.585 143.005 ;
        RECT 1034.705 142.995 1035.085 143.030 ;
        RECT 1037.750 142.995 1039.085 143.375 ;
        RECT 1042.705 143.355 1043.085 143.375 ;
        RECT 1040.240 143.035 1043.150 143.355 ;
        RECT 1059.640 143.250 1060.020 143.285 ;
        RECT 1042.705 142.995 1043.085 143.035 ;
        RECT 1059.375 142.940 1062.385 143.250 ;
        RECT 1059.640 142.905 1060.020 142.940 ;
        RECT 1063.640 142.905 1064.730 143.285 ;
        RECT 1067.640 143.280 1068.020 143.285 ;
        RECT 1065.160 142.915 1068.025 143.280 ;
        RECT 1073.140 143.260 1073.520 143.285 ;
        RECT 1073.125 142.940 1075.270 143.260 ;
        RECT 1067.640 142.905 1068.020 142.915 ;
        RECT 1073.140 142.905 1073.520 142.940 ;
        RECT 1076.185 142.905 1077.520 143.285 ;
        RECT 1081.140 143.265 1081.520 143.285 ;
        RECT 1078.675 142.945 1081.585 143.265 ;
        RECT 1081.140 142.905 1081.520 142.945 ;
        RECT 1085.770 142.765 1086.150 143.145 ;
        RECT 1088.175 142.780 1089.955 143.070 ;
        RECT 1091.430 142.870 1092.620 143.155 ;
        RECT 1095.550 142.750 1096.860 143.070 ;
        RECT 1004.375 142.255 1004.755 142.635 ;
        RECT 1008.120 142.295 1008.500 142.675 ;
        RECT 1010.830 142.285 1011.210 142.665 ;
        RECT 1012.240 142.130 1015.420 142.450 ;
        RECT 1086.905 142.165 1087.285 142.545 ;
        RECT 1090.650 142.205 1091.030 142.585 ;
        RECT 1093.360 142.195 1093.740 142.575 ;
        RECT 1019.555 141.685 1021.045 142.065 ;
        RECT 1021.745 141.685 1023.030 142.065 ;
        RECT 1041.060 141.685 1042.545 142.065 ;
        RECT 1043.245 141.685 1044.320 142.065 ;
        RECT 1094.770 142.040 1097.950 142.360 ;
        RECT 1057.990 141.595 1059.480 141.975 ;
        RECT 1081.680 141.595 1082.755 141.975 ;
        RECT 1021.205 140.995 1022.295 141.375 ;
        RECT 1023.250 141.005 1024.770 141.365 ;
        RECT 1025.690 141.000 1038.540 141.335 ;
        RECT 1042.705 141.330 1043.085 141.375 ;
        RECT 1041.970 141.030 1043.280 141.330 ;
        RECT 1042.705 140.995 1043.085 141.030 ;
        RECT 1059.640 140.905 1060.730 141.285 ;
        RECT 1061.685 140.915 1063.205 141.275 ;
        RECT 1064.125 140.910 1076.975 141.245 ;
        RECT 1081.140 141.240 1081.520 141.285 ;
        RECT 1080.405 140.940 1081.715 141.240 ;
        RECT 1081.140 140.905 1081.520 140.940 ;
        RECT 1018.060 140.410 1051.140 140.485 ;
        RECT 1018.060 140.135 1083.150 140.410 ;
        RECT 1050.200 140.045 1083.150 140.135 ;
        RECT 1084.945 140.035 1089.205 140.390 ;
        RECT 1002.170 139.540 1006.265 139.545 ;
        RECT 985.590 139.535 990.805 139.540 ;
        RECT 1001.050 139.535 1006.265 139.540 ;
        RECT 1016.510 139.535 1056.760 139.540 ;
        RECT 985.590 139.450 1056.760 139.535 ;
        RECT 1083.150 139.450 1088.795 139.455 ;
        RECT 1099.410 139.450 1099.790 145.280 ;
        RECT 1108.290 145.230 1112.790 145.540 ;
        RECT 1184.675 145.370 1188.805 145.670 ;
        RECT 1104.250 144.680 1110.640 144.970 ;
        RECT 1103.665 144.100 1119.685 144.435 ;
        RECT 1168.595 144.350 1174.510 144.685 ;
        RECT 1171.865 144.330 1174.510 144.350 ;
        RECT 1103.015 143.515 1105.935 143.815 ;
        RECT 1109.480 143.500 1112.850 143.800 ;
        RECT 1149.190 143.710 1152.490 144.090 ;
        RECT 1153.190 143.710 1156.490 144.090 ;
        RECT 1162.690 143.710 1165.990 144.090 ;
        RECT 1166.690 143.710 1169.990 144.090 ;
        RECT 1101.230 142.765 1101.610 143.145 ;
        RECT 1103.635 142.780 1105.415 143.070 ;
        RECT 1106.890 142.870 1108.080 143.155 ;
        RECT 1111.010 142.750 1112.320 143.070 ;
        RECT 1102.365 142.165 1102.745 142.545 ;
        RECT 1106.110 142.205 1106.490 142.585 ;
        RECT 1108.820 142.195 1109.200 142.575 ;
        RECT 1110.230 142.040 1113.410 142.360 ;
        RECT 1149.190 141.710 1150.475 142.090 ;
        RECT 1168.505 141.710 1169.990 142.090 ;
        RECT 1100.510 140.955 1104.660 141.225 ;
        RECT 1150.695 141.030 1152.215 141.390 ;
        RECT 1100.160 139.450 1104.255 139.455 ;
        RECT 985.590 139.445 1088.795 139.450 ;
        RECT 1099.040 139.445 1104.255 139.450 ;
        RECT 985.590 138.640 1114.070 139.445 ;
        RECT 1145.505 138.665 1172.160 139.565 ;
        RECT 1182.300 139.540 1182.680 145.370 ;
        RECT 1191.180 145.320 1195.680 145.630 ;
        RECT 1200.135 145.370 1204.265 145.670 ;
        RECT 1187.140 144.770 1193.530 145.060 ;
        RECT 1186.555 144.190 1197.210 144.525 ;
        RECT 1185.905 143.605 1188.825 143.905 ;
        RECT 1192.370 143.590 1195.740 143.890 ;
        RECT 1184.120 142.855 1184.500 143.235 ;
        RECT 1186.525 142.870 1188.305 143.160 ;
        RECT 1189.780 142.960 1190.970 143.245 ;
        RECT 1193.900 142.840 1195.210 143.160 ;
        RECT 1185.255 142.255 1185.635 142.635 ;
        RECT 1189.000 142.295 1189.380 142.675 ;
        RECT 1191.710 142.285 1192.090 142.665 ;
        RECT 1193.120 142.130 1196.300 142.450 ;
        RECT 1183.050 139.540 1187.145 139.545 ;
        RECT 1197.760 139.540 1198.140 145.370 ;
        RECT 1206.640 145.320 1211.140 145.630 ;
        RECT 1282.665 145.280 1286.795 145.580 ;
        RECT 1289.170 145.230 1293.670 145.540 ;
        RECT 1298.125 145.280 1302.255 145.580 ;
        RECT 1213.870 145.070 1249.780 145.160 ;
        RECT 1202.600 144.770 1208.990 145.060 ;
        RECT 1213.870 144.890 1280.910 145.070 ;
        RECT 1249.165 144.800 1280.910 144.890 ;
        RECT 1285.130 144.680 1291.520 144.970 ;
        RECT 1202.015 144.190 1212.520 144.525 ;
        RECT 1237.490 144.325 1248.040 144.660 ;
        RECT 1275.925 144.235 1279.870 144.570 ;
        RECT 1284.545 144.100 1295.025 144.435 ;
        RECT 1201.365 143.605 1204.285 143.905 ;
        RECT 1207.830 143.590 1211.200 143.890 ;
        RECT 1216.080 143.685 1217.385 144.065 ;
        RECT 1218.085 143.685 1221.385 144.065 ;
        RECT 1222.085 143.685 1225.385 144.065 ;
        RECT 1226.085 143.685 1227.445 144.065 ;
        RECT 1229.420 143.685 1230.885 144.065 ;
        RECT 1231.585 143.685 1234.885 144.065 ;
        RECT 1235.585 143.685 1238.885 144.065 ;
        RECT 1239.585 143.685 1240.765 144.065 ;
        RECT 1254.515 143.595 1255.820 143.975 ;
        RECT 1256.520 143.595 1259.820 143.975 ;
        RECT 1260.520 143.595 1263.820 143.975 ;
        RECT 1264.520 143.595 1265.880 143.975 ;
        RECT 1267.855 143.595 1269.320 143.975 ;
        RECT 1270.020 143.595 1273.320 143.975 ;
        RECT 1274.020 143.595 1277.320 143.975 ;
        RECT 1278.020 143.595 1279.200 143.975 ;
        RECT 1283.895 143.515 1286.815 143.815 ;
        RECT 1290.360 143.500 1293.730 143.800 ;
        RECT 1217.545 143.340 1217.925 143.375 ;
        RECT 1199.580 142.855 1199.960 143.235 ;
        RECT 1201.985 142.870 1203.765 143.160 ;
        RECT 1205.240 142.960 1206.430 143.245 ;
        RECT 1209.360 142.840 1210.670 143.160 ;
        RECT 1217.280 143.030 1220.290 143.340 ;
        RECT 1217.545 142.995 1217.925 143.030 ;
        RECT 1221.545 142.995 1222.635 143.375 ;
        RECT 1225.545 143.370 1225.925 143.375 ;
        RECT 1223.065 143.005 1225.930 143.370 ;
        RECT 1231.045 143.350 1231.425 143.375 ;
        RECT 1231.030 143.030 1233.175 143.350 ;
        RECT 1225.545 142.995 1225.925 143.005 ;
        RECT 1231.045 142.995 1231.425 143.030 ;
        RECT 1234.090 142.995 1235.425 143.375 ;
        RECT 1239.045 143.355 1239.425 143.375 ;
        RECT 1236.580 143.035 1239.490 143.355 ;
        RECT 1255.980 143.250 1256.360 143.285 ;
        RECT 1239.045 142.995 1239.425 143.035 ;
        RECT 1255.715 142.940 1258.725 143.250 ;
        RECT 1255.980 142.905 1256.360 142.940 ;
        RECT 1259.980 142.905 1261.070 143.285 ;
        RECT 1263.980 143.280 1264.360 143.285 ;
        RECT 1261.500 142.915 1264.365 143.280 ;
        RECT 1269.480 143.260 1269.860 143.285 ;
        RECT 1269.465 142.940 1271.610 143.260 ;
        RECT 1263.980 142.905 1264.360 142.915 ;
        RECT 1269.480 142.905 1269.860 142.940 ;
        RECT 1272.525 142.905 1273.860 143.285 ;
        RECT 1277.480 143.265 1277.860 143.285 ;
        RECT 1275.015 142.945 1277.925 143.265 ;
        RECT 1277.480 142.905 1277.860 142.945 ;
        RECT 1282.110 142.765 1282.490 143.145 ;
        RECT 1284.515 142.780 1286.295 143.070 ;
        RECT 1287.770 142.870 1288.960 143.155 ;
        RECT 1291.890 142.750 1293.200 143.070 ;
        RECT 1200.715 142.255 1201.095 142.635 ;
        RECT 1204.460 142.295 1204.840 142.675 ;
        RECT 1207.170 142.285 1207.550 142.665 ;
        RECT 1208.580 142.130 1211.760 142.450 ;
        RECT 1283.245 142.165 1283.625 142.545 ;
        RECT 1286.990 142.205 1287.370 142.585 ;
        RECT 1289.700 142.195 1290.080 142.575 ;
        RECT 1215.895 141.685 1217.385 142.065 ;
        RECT 1218.085 141.685 1219.370 142.065 ;
        RECT 1237.400 141.685 1238.885 142.065 ;
        RECT 1239.585 141.685 1240.660 142.065 ;
        RECT 1291.110 142.040 1294.290 142.360 ;
        RECT 1254.330 141.595 1255.820 141.975 ;
        RECT 1256.520 141.595 1257.805 141.975 ;
        RECT 1275.835 141.595 1277.320 141.975 ;
        RECT 1278.020 141.595 1279.095 141.975 ;
        RECT 1217.545 140.995 1218.635 141.375 ;
        RECT 1219.590 141.005 1221.110 141.365 ;
        RECT 1222.030 141.000 1234.880 141.335 ;
        RECT 1239.045 141.330 1239.425 141.375 ;
        RECT 1238.310 141.030 1239.620 141.330 ;
        RECT 1239.045 140.995 1239.425 141.030 ;
        RECT 1255.980 140.905 1257.070 141.285 ;
        RECT 1258.025 140.915 1259.545 141.275 ;
        RECT 1260.465 140.910 1273.315 141.245 ;
        RECT 1277.480 141.240 1277.860 141.285 ;
        RECT 1276.745 140.940 1278.055 141.240 ;
        RECT 1277.480 140.905 1277.860 140.940 ;
        RECT 1214.400 140.410 1247.480 140.485 ;
        RECT 1214.400 140.135 1279.490 140.410 ;
        RECT 1246.540 140.045 1279.490 140.135 ;
        RECT 1281.285 140.035 1285.545 140.390 ;
        RECT 1198.510 139.540 1202.605 139.545 ;
        RECT 1181.930 139.535 1187.145 139.540 ;
        RECT 1197.390 139.535 1202.605 139.540 ;
        RECT 1212.850 139.535 1253.100 139.540 ;
        RECT 1181.930 139.450 1253.100 139.535 ;
        RECT 1279.490 139.450 1285.135 139.455 ;
        RECT 1295.750 139.450 1296.130 145.280 ;
        RECT 1304.630 145.230 1309.130 145.540 ;
        RECT 1300.590 144.680 1306.980 144.970 ;
        RECT 1299.355 143.515 1302.275 143.815 ;
        RECT 1305.820 143.500 1309.190 143.800 ;
        RECT 1297.570 142.765 1297.950 143.145 ;
        RECT 1303.230 142.870 1304.420 143.155 ;
        RECT 1302.450 142.205 1302.830 142.585 ;
        RECT 1306.570 142.040 1309.750 142.360 ;
        RECT 1296.850 140.955 1301.000 141.225 ;
        RECT 1296.500 139.450 1300.595 139.455 ;
        RECT 1181.930 139.445 1285.135 139.450 ;
        RECT 1295.380 139.445 1300.595 139.450 ;
        RECT 1181.930 138.640 1310.410 139.445 ;
        RECT 467.440 138.515 525.015 138.605 ;
        RECT 663.815 138.550 721.390 138.640 ;
        RECT 860.155 138.550 917.730 138.640 ;
        RECT 1056.495 138.550 1114.070 138.640 ;
        RECT 1252.835 138.550 1310.410 138.640 ;
        RECT 3.960 134.845 76.350 134.870 ;
        RECT 200.325 134.845 272.715 134.870 ;
        RECT -81.495 133.795 -56.060 134.695 ;
        RECT -31.170 133.875 -5.735 134.775 ;
        RECT 3.960 133.970 132.405 134.845 ;
        RECT -79.010 131.615 -77.810 131.995 ;
        RECT -76.055 131.400 -73.780 131.910 ;
        RECT -71.155 131.400 -68.855 131.910 ;
        RECT -66.560 131.400 -64.280 131.910 ;
        RECT -59.485 131.715 -58.250 132.095 ;
        RECT -28.685 131.695 -27.485 132.075 ;
        RECT -25.730 131.480 -23.455 131.990 ;
        RECT -20.830 131.480 -18.530 131.990 ;
        RECT -16.235 131.480 -13.955 131.990 ;
        RECT -9.160 131.795 -7.925 132.175 ;
        RECT -79.010 129.315 -75.750 129.695 ;
        RECT -75.010 129.315 -71.750 129.695 ;
        RECT -65.510 129.315 -62.250 129.695 ;
        RECT -61.510 129.315 -58.250 129.695 ;
        RECT -28.685 129.395 -25.425 129.775 ;
        RECT -24.685 129.395 -21.425 129.775 ;
        RECT -15.185 129.395 -11.925 129.775 ;
        RECT -11.185 129.395 -7.925 129.775 ;
        RECT -78.345 127.730 -56.060 127.740 ;
        RECT -78.345 127.400 -54.520 127.730 ;
        RECT -28.020 127.480 -1.725 127.820 ;
        RECT -56.280 127.380 -54.520 127.400 ;
        RECT 4.330 126.810 4.710 133.970 ;
        RECT 6.160 129.755 9.535 130.155 ;
        RECT 9.905 129.515 10.285 129.895 ;
        RECT 12.620 129.555 13.000 129.935 ;
        RECT 16.805 129.505 17.185 129.885 ;
        RECT 7.230 129.090 8.970 129.380 ;
        RECT 11.020 129.040 12.220 129.330 ;
        RECT 13.730 129.010 16.340 129.435 ;
        RECT 17.940 129.105 18.320 129.485 ;
        RECT 5.475 128.330 19.040 128.645 ;
        RECT 5.470 127.585 19.030 127.885 ;
        RECT 5.490 126.870 12.215 127.170 ;
        RECT 15.915 126.570 19.020 126.845 ;
        RECT 19.790 126.810 20.170 133.970 ;
        RECT 76.050 133.945 132.405 133.970 ;
        RECT 36.430 132.960 73.980 132.985 ;
        RECT 36.430 132.700 101.810 132.960 ;
        RECT 73.035 132.675 101.810 132.700 ;
        RECT 103.480 132.655 110.185 132.955 ;
        RECT 37.940 131.790 39.395 132.170 ;
        RECT 40.135 131.790 41.335 132.170 ;
        RECT 43.090 131.575 45.365 132.085 ;
        RECT 47.990 131.575 50.290 132.085 ;
        RECT 52.585 131.575 54.865 132.085 ;
        RECT 59.660 131.890 60.895 132.270 ;
        RECT 61.635 131.890 62.915 132.270 ;
        RECT 76.340 131.765 77.795 132.145 ;
        RECT 61.075 131.535 61.455 131.570 ;
        RECT 81.490 131.550 83.765 132.060 ;
        RECT 86.390 131.550 88.690 132.060 ;
        RECT 90.985 131.550 93.265 132.060 ;
        RECT 100.035 131.865 101.315 132.245 ;
        RECT 39.575 131.430 39.955 131.470 ;
        RECT 39.505 131.125 42.340 131.430 ;
        RECT 58.320 131.225 61.455 131.535 ;
        RECT 99.475 131.510 99.855 131.545 ;
        RECT 77.975 131.405 78.355 131.445 ;
        RECT 61.075 131.190 61.455 131.225 ;
        RECT 39.575 131.090 39.955 131.125 ;
        RECT 77.905 131.100 80.740 131.405 ;
        RECT 96.720 131.200 99.855 131.510 ;
        RECT 99.475 131.165 99.855 131.200 ;
        RECT 77.975 131.065 78.355 131.100 ;
        RECT 21.620 129.715 25.025 130.155 ;
        RECT 25.365 129.515 25.745 129.895 ;
        RECT 28.080 129.555 28.460 129.935 ;
        RECT 32.265 129.505 32.645 129.885 ;
        RECT 38.100 129.490 39.395 129.870 ;
        RECT 40.135 129.490 43.395 129.870 ;
        RECT 44.135 129.490 47.395 129.870 ;
        RECT 48.135 129.490 49.320 129.870 ;
        RECT 51.585 129.490 52.895 129.870 ;
        RECT 53.635 129.490 56.895 129.870 ;
        RECT 57.635 129.490 60.895 129.870 ;
        RECT 61.635 129.490 62.650 129.870 ;
        RECT 22.690 129.090 24.430 129.380 ;
        RECT 26.480 129.040 27.680 129.330 ;
        RECT 29.190 129.010 31.785 129.385 ;
        RECT 33.400 129.105 33.780 129.485 ;
        RECT 76.500 129.465 77.795 129.845 ;
        RECT 82.535 129.465 85.795 129.845 ;
        RECT 86.535 129.465 87.720 129.845 ;
        RECT 89.985 129.465 91.295 129.845 ;
        RECT 92.035 129.465 95.295 129.845 ;
        RECT 100.035 129.465 101.050 129.845 ;
        RECT 104.115 129.710 107.530 130.130 ;
        RECT 107.860 129.490 108.240 129.870 ;
        RECT 110.575 129.530 110.955 129.910 ;
        RECT 114.760 129.480 115.140 129.860 ;
        RECT 39.575 128.790 39.955 129.170 ;
        RECT 43.575 128.790 43.955 129.170 ;
        RECT 47.575 129.125 47.955 129.170 ;
        RECT 53.075 129.125 53.455 129.170 ;
        RECT 47.525 128.810 53.460 129.125 ;
        RECT 47.575 128.790 47.955 128.810 ;
        RECT 53.075 128.790 53.455 128.810 ;
        RECT 57.075 128.790 57.455 129.170 ;
        RECT 61.075 128.790 61.455 129.170 ;
        RECT 77.975 128.765 78.355 129.145 ;
        RECT 81.975 128.765 82.355 129.145 ;
        RECT 85.975 129.100 86.355 129.145 ;
        RECT 91.475 129.100 91.855 129.145 ;
        RECT 85.925 128.785 91.860 129.100 ;
        RECT 85.975 128.765 86.355 128.785 ;
        RECT 91.475 128.765 91.855 128.785 ;
        RECT 95.475 128.765 95.855 129.145 ;
        RECT 99.475 128.765 99.855 129.145 ;
        RECT 105.185 129.065 106.925 129.355 ;
        RECT 108.975 129.015 110.175 129.305 ;
        RECT 111.685 128.975 114.315 129.430 ;
        RECT 115.895 129.080 116.275 129.460 ;
        RECT 20.930 128.330 34.755 128.630 ;
        RECT 36.430 128.165 52.440 128.540 ;
        RECT 70.065 128.140 90.840 128.515 ;
        RECT 20.935 127.585 39.355 127.885 ;
        RECT 40.800 127.575 68.110 127.915 ;
        RECT 20.415 126.870 27.675 127.170 ;
        RECT 5.470 126.250 9.595 126.520 ;
        RECT 20.970 126.335 25.055 126.605 ;
        RECT 31.375 126.570 35.125 126.845 ;
        RECT 36.430 126.810 62.660 127.200 ;
        RECT 69.095 126.785 101.060 127.175 ;
        RECT 113.870 126.545 117.000 126.820 ;
        RECT 117.745 126.785 118.125 133.945 ;
        RECT 165.000 133.885 190.435 134.785 ;
        RECT 200.325 133.970 328.770 134.845 ;
        RECT 593.100 134.830 665.490 134.855 ;
        RECT 789.440 134.830 861.830 134.855 ;
        RECT 985.780 134.830 1058.170 134.855 ;
        RECT 1182.120 134.830 1254.510 134.855 ;
        RECT 396.725 134.795 469.115 134.820 ;
        RECT 118.985 131.485 125.725 131.785 ;
        RECT 167.485 131.705 168.685 132.085 ;
        RECT 170.440 131.490 172.715 132.000 ;
        RECT 175.340 131.490 177.640 132.000 ;
        RECT 179.935 131.490 182.215 132.000 ;
        RECT 187.010 131.805 188.245 132.185 ;
        RECT 119.575 129.690 123.030 130.130 ;
        RECT 123.320 129.490 123.700 129.870 ;
        RECT 126.035 129.530 126.415 129.910 ;
        RECT 130.220 129.480 130.600 129.860 ;
        RECT 120.645 129.065 122.385 129.355 ;
        RECT 124.435 129.015 125.635 129.305 ;
        RECT 127.145 128.985 129.770 129.395 ;
        RECT 131.355 129.080 131.735 129.460 ;
        RECT 167.485 129.405 170.745 129.785 ;
        RECT 171.485 129.405 174.745 129.785 ;
        RECT 180.985 129.405 184.245 129.785 ;
        RECT 184.985 129.405 188.245 129.785 ;
        RECT 118.390 128.305 134.310 128.605 ;
        RECT 118.925 127.560 135.870 127.860 ;
        RECT 168.150 127.490 194.445 127.830 ;
        RECT 129.330 126.545 137.030 126.820 ;
        RECT 200.695 126.810 201.075 133.970 ;
        RECT 202.525 129.755 205.900 130.155 ;
        RECT 206.270 129.515 206.650 129.895 ;
        RECT 208.985 129.555 209.365 129.935 ;
        RECT 213.170 129.505 213.550 129.885 ;
        RECT 203.595 129.090 205.335 129.380 ;
        RECT 207.385 129.040 208.585 129.330 ;
        RECT 210.095 129.010 212.705 129.435 ;
        RECT 214.305 129.105 214.685 129.485 ;
        RECT 201.840 128.330 215.405 128.645 ;
        RECT 201.835 127.585 215.395 127.885 ;
        RECT 201.855 126.870 208.580 127.170 ;
        RECT 212.280 126.570 215.385 126.845 ;
        RECT 216.155 126.810 216.535 133.970 ;
        RECT 272.415 133.945 328.770 133.970 ;
        RECT 232.795 132.960 270.345 132.985 ;
        RECT 232.795 132.700 298.175 132.960 ;
        RECT 269.400 132.675 298.175 132.700 ;
        RECT 299.845 132.655 306.550 132.955 ;
        RECT 234.305 131.790 235.760 132.170 ;
        RECT 236.500 131.790 237.700 132.170 ;
        RECT 239.455 131.575 241.730 132.085 ;
        RECT 244.355 131.575 246.655 132.085 ;
        RECT 248.950 131.575 251.230 132.085 ;
        RECT 256.025 131.890 257.260 132.270 ;
        RECT 258.000 131.890 259.280 132.270 ;
        RECT 272.705 131.765 274.160 132.145 ;
        RECT 257.440 131.535 257.820 131.570 ;
        RECT 277.855 131.550 280.130 132.060 ;
        RECT 282.755 131.550 285.055 132.060 ;
        RECT 287.350 131.550 289.630 132.060 ;
        RECT 296.400 131.865 297.680 132.245 ;
        RECT 235.940 131.430 236.320 131.470 ;
        RECT 235.870 131.125 238.705 131.430 ;
        RECT 254.685 131.225 257.820 131.535 ;
        RECT 295.840 131.510 296.220 131.545 ;
        RECT 274.340 131.405 274.720 131.445 ;
        RECT 257.440 131.190 257.820 131.225 ;
        RECT 235.940 131.090 236.320 131.125 ;
        RECT 274.270 131.100 277.105 131.405 ;
        RECT 293.085 131.200 296.220 131.510 ;
        RECT 295.840 131.165 296.220 131.200 ;
        RECT 274.340 131.065 274.720 131.100 ;
        RECT 217.985 129.715 221.390 130.155 ;
        RECT 221.730 129.515 222.110 129.895 ;
        RECT 224.445 129.555 224.825 129.935 ;
        RECT 228.630 129.505 229.010 129.885 ;
        RECT 234.465 129.490 235.760 129.870 ;
        RECT 236.500 129.490 239.760 129.870 ;
        RECT 240.500 129.490 243.760 129.870 ;
        RECT 244.500 129.490 245.685 129.870 ;
        RECT 247.950 129.490 249.260 129.870 ;
        RECT 250.000 129.490 253.260 129.870 ;
        RECT 254.000 129.490 257.260 129.870 ;
        RECT 258.000 129.490 259.015 129.870 ;
        RECT 219.055 129.090 220.795 129.380 ;
        RECT 222.845 129.040 224.045 129.330 ;
        RECT 225.555 129.010 228.150 129.385 ;
        RECT 229.765 129.105 230.145 129.485 ;
        RECT 272.865 129.465 274.160 129.845 ;
        RECT 278.900 129.465 282.160 129.845 ;
        RECT 282.900 129.465 284.085 129.845 ;
        RECT 286.350 129.465 287.660 129.845 ;
        RECT 288.400 129.465 291.660 129.845 ;
        RECT 296.400 129.465 297.415 129.845 ;
        RECT 300.480 129.710 303.895 130.130 ;
        RECT 304.225 129.490 304.605 129.870 ;
        RECT 306.940 129.530 307.320 129.910 ;
        RECT 311.125 129.480 311.505 129.860 ;
        RECT 235.940 128.790 236.320 129.170 ;
        RECT 239.940 128.790 240.320 129.170 ;
        RECT 243.940 129.125 244.320 129.170 ;
        RECT 249.440 129.125 249.820 129.170 ;
        RECT 243.890 128.810 249.825 129.125 ;
        RECT 243.940 128.790 244.320 128.810 ;
        RECT 249.440 128.790 249.820 128.810 ;
        RECT 253.440 128.790 253.820 129.170 ;
        RECT 257.440 128.790 257.820 129.170 ;
        RECT 274.340 128.765 274.720 129.145 ;
        RECT 278.340 128.765 278.720 129.145 ;
        RECT 282.340 129.100 282.720 129.145 ;
        RECT 287.840 129.100 288.220 129.145 ;
        RECT 282.290 128.785 288.225 129.100 ;
        RECT 282.340 128.765 282.720 128.785 ;
        RECT 287.840 128.765 288.220 128.785 ;
        RECT 291.840 128.765 292.220 129.145 ;
        RECT 295.840 128.765 296.220 129.145 ;
        RECT 301.550 129.065 303.290 129.355 ;
        RECT 305.340 129.015 306.540 129.305 ;
        RECT 308.050 128.975 310.680 129.430 ;
        RECT 312.260 129.080 312.640 129.460 ;
        RECT 217.295 128.330 231.120 128.630 ;
        RECT 232.795 128.165 248.805 128.540 ;
        RECT 266.430 128.140 287.205 128.515 ;
        RECT 217.300 127.585 235.720 127.885 ;
        RECT 237.165 127.575 264.475 127.915 ;
        RECT 216.780 126.870 224.040 127.170 ;
        RECT 36.430 126.445 55.100 126.455 ;
        RECT 36.430 126.430 66.450 126.445 ;
        RECT 36.430 126.420 93.500 126.430 ;
        RECT 36.430 126.135 102.505 126.420 ;
        RECT 201.835 126.250 205.960 126.520 ;
        RECT 217.335 126.335 221.420 126.605 ;
        RECT 227.740 126.570 231.490 126.845 ;
        RECT 232.795 126.810 259.025 127.200 ;
        RECT 265.460 126.785 297.425 127.175 ;
        RECT 310.235 126.545 313.365 126.820 ;
        RECT 314.110 126.785 314.490 133.945 ;
        RECT 361.390 133.845 386.825 134.745 ;
        RECT 396.725 133.920 525.170 134.795 ;
        RECT 315.350 131.485 322.090 131.785 ;
        RECT 363.875 131.665 365.075 132.045 ;
        RECT 366.830 131.450 369.105 131.960 ;
        RECT 371.730 131.450 374.030 131.960 ;
        RECT 376.325 131.450 378.605 131.960 ;
        RECT 383.400 131.765 384.635 132.145 ;
        RECT 315.940 129.690 319.395 130.130 ;
        RECT 319.685 129.490 320.065 129.870 ;
        RECT 322.400 129.530 322.780 129.910 ;
        RECT 326.585 129.480 326.965 129.860 ;
        RECT 317.010 129.065 318.750 129.355 ;
        RECT 320.800 129.015 322.000 129.305 ;
        RECT 323.510 128.985 326.135 129.395 ;
        RECT 327.720 129.080 328.100 129.460 ;
        RECT 363.875 129.365 367.135 129.745 ;
        RECT 367.875 129.365 371.135 129.745 ;
        RECT 377.375 129.365 380.635 129.745 ;
        RECT 381.375 129.365 384.635 129.745 ;
        RECT 314.755 128.305 330.675 128.605 ;
        RECT 315.290 127.560 332.235 127.860 ;
        RECT 364.540 127.450 390.835 127.790 ;
        RECT 325.695 126.545 333.395 126.820 ;
        RECT 397.095 126.760 397.475 133.920 ;
        RECT 398.925 129.705 402.300 130.105 ;
        RECT 402.670 129.465 403.050 129.845 ;
        RECT 405.385 129.505 405.765 129.885 ;
        RECT 409.570 129.455 409.950 129.835 ;
        RECT 399.995 129.040 401.735 129.330 ;
        RECT 403.785 128.990 404.985 129.280 ;
        RECT 406.495 128.960 409.105 129.385 ;
        RECT 410.705 129.055 411.085 129.435 ;
        RECT 398.240 128.280 411.805 128.595 ;
        RECT 398.235 127.535 411.795 127.835 ;
        RECT 398.255 126.820 404.980 127.120 ;
        RECT 408.680 126.520 411.785 126.795 ;
        RECT 412.555 126.760 412.935 133.920 ;
        RECT 468.815 133.895 525.170 133.920 ;
        RECT 429.195 132.910 466.745 132.935 ;
        RECT 429.195 132.650 494.575 132.910 ;
        RECT 465.800 132.625 494.575 132.650 ;
        RECT 496.245 132.605 502.950 132.905 ;
        RECT 430.705 131.740 432.160 132.120 ;
        RECT 432.900 131.740 434.100 132.120 ;
        RECT 435.855 131.525 438.130 132.035 ;
        RECT 440.755 131.525 443.055 132.035 ;
        RECT 445.350 131.525 447.630 132.035 ;
        RECT 452.425 131.840 453.660 132.220 ;
        RECT 454.400 131.840 455.680 132.220 ;
        RECT 469.105 131.715 470.560 132.095 ;
        RECT 453.840 131.485 454.220 131.520 ;
        RECT 474.255 131.500 476.530 132.010 ;
        RECT 479.155 131.500 481.455 132.010 ;
        RECT 483.750 131.500 486.030 132.010 ;
        RECT 492.800 131.815 494.080 132.195 ;
        RECT 432.340 131.380 432.720 131.420 ;
        RECT 432.270 131.075 435.105 131.380 ;
        RECT 451.085 131.175 454.220 131.485 ;
        RECT 492.240 131.460 492.620 131.495 ;
        RECT 470.740 131.355 471.120 131.395 ;
        RECT 453.840 131.140 454.220 131.175 ;
        RECT 432.340 131.040 432.720 131.075 ;
        RECT 470.670 131.050 473.505 131.355 ;
        RECT 489.485 131.150 492.620 131.460 ;
        RECT 492.240 131.115 492.620 131.150 ;
        RECT 470.740 131.015 471.120 131.050 ;
        RECT 414.385 129.665 417.790 130.105 ;
        RECT 418.130 129.465 418.510 129.845 ;
        RECT 420.845 129.505 421.225 129.885 ;
        RECT 425.030 129.455 425.410 129.835 ;
        RECT 430.865 129.440 432.160 129.820 ;
        RECT 432.900 129.440 436.160 129.820 ;
        RECT 436.900 129.440 440.160 129.820 ;
        RECT 440.900 129.440 442.085 129.820 ;
        RECT 444.350 129.440 445.660 129.820 ;
        RECT 446.400 129.440 449.660 129.820 ;
        RECT 450.400 129.440 453.660 129.820 ;
        RECT 454.400 129.440 455.415 129.820 ;
        RECT 415.455 129.040 417.195 129.330 ;
        RECT 419.245 128.990 420.445 129.280 ;
        RECT 421.955 128.960 424.550 129.335 ;
        RECT 426.165 129.055 426.545 129.435 ;
        RECT 469.265 129.415 470.560 129.795 ;
        RECT 475.300 129.415 478.560 129.795 ;
        RECT 479.300 129.415 480.485 129.795 ;
        RECT 482.750 129.415 484.060 129.795 ;
        RECT 484.800 129.415 488.060 129.795 ;
        RECT 492.800 129.415 493.815 129.795 ;
        RECT 496.880 129.660 500.295 130.080 ;
        RECT 500.625 129.440 501.005 129.820 ;
        RECT 503.340 129.480 503.720 129.860 ;
        RECT 507.525 129.430 507.905 129.810 ;
        RECT 432.340 128.740 432.720 129.120 ;
        RECT 436.340 128.740 436.720 129.120 ;
        RECT 440.340 129.075 440.720 129.120 ;
        RECT 445.840 129.075 446.220 129.120 ;
        RECT 440.290 128.760 446.225 129.075 ;
        RECT 440.340 128.740 440.720 128.760 ;
        RECT 445.840 128.740 446.220 128.760 ;
        RECT 449.840 128.740 450.220 129.120 ;
        RECT 453.840 128.740 454.220 129.120 ;
        RECT 470.740 128.715 471.120 129.095 ;
        RECT 474.740 128.715 475.120 129.095 ;
        RECT 478.740 129.050 479.120 129.095 ;
        RECT 484.240 129.050 484.620 129.095 ;
        RECT 478.690 128.735 484.625 129.050 ;
        RECT 478.740 128.715 479.120 128.735 ;
        RECT 484.240 128.715 484.620 128.735 ;
        RECT 488.240 128.715 488.620 129.095 ;
        RECT 492.240 128.715 492.620 129.095 ;
        RECT 497.950 129.015 499.690 129.305 ;
        RECT 501.740 128.965 502.940 129.255 ;
        RECT 504.450 128.925 507.080 129.380 ;
        RECT 508.660 129.030 509.040 129.410 ;
        RECT 413.695 128.280 427.520 128.580 ;
        RECT 429.195 128.115 445.205 128.490 ;
        RECT 462.830 128.090 483.605 128.465 ;
        RECT 413.700 127.535 432.120 127.835 ;
        RECT 433.565 127.525 460.875 127.865 ;
        RECT 413.180 126.820 420.440 127.120 ;
        RECT 232.795 126.445 251.465 126.455 ;
        RECT 232.795 126.430 262.815 126.445 ;
        RECT 232.795 126.420 289.865 126.430 ;
        RECT 232.795 126.135 298.870 126.420 ;
        RECT 398.235 126.200 402.360 126.470 ;
        RECT 413.735 126.285 417.820 126.555 ;
        RECT 424.140 126.520 427.890 126.795 ;
        RECT 429.195 126.760 455.425 127.150 ;
        RECT 461.860 126.735 493.825 127.125 ;
        RECT 506.635 126.495 509.765 126.770 ;
        RECT 510.510 126.735 510.890 133.895 ;
        RECT 557.710 133.890 583.145 134.790 ;
        RECT 593.100 133.955 721.545 134.830 ;
        RECT 511.750 131.435 518.490 131.735 ;
        RECT 560.195 131.710 561.395 132.090 ;
        RECT 563.150 131.495 565.425 132.005 ;
        RECT 568.050 131.495 570.350 132.005 ;
        RECT 572.645 131.495 574.925 132.005 ;
        RECT 579.720 131.810 580.955 132.190 ;
        RECT 512.340 129.640 515.795 130.080 ;
        RECT 516.085 129.440 516.465 129.820 ;
        RECT 518.800 129.480 519.180 129.860 ;
        RECT 522.985 129.430 523.365 129.810 ;
        RECT 560.195 129.410 563.455 129.790 ;
        RECT 564.195 129.410 567.455 129.790 ;
        RECT 573.695 129.410 576.955 129.790 ;
        RECT 577.695 129.410 580.955 129.790 ;
        RECT 513.410 129.015 515.150 129.305 ;
        RECT 517.200 128.965 518.400 129.255 ;
        RECT 519.910 128.935 522.535 129.345 ;
        RECT 524.120 129.030 524.500 129.410 ;
        RECT 511.155 128.255 527.075 128.555 ;
        RECT 511.690 127.510 528.635 127.810 ;
        RECT 560.860 127.495 587.155 127.835 ;
        RECT 593.470 126.795 593.850 133.955 ;
        RECT 595.300 129.740 598.675 130.140 ;
        RECT 599.045 129.500 599.425 129.880 ;
        RECT 601.760 129.540 602.140 129.920 ;
        RECT 605.945 129.490 606.325 129.870 ;
        RECT 596.370 129.075 598.110 129.365 ;
        RECT 600.160 129.025 601.360 129.315 ;
        RECT 602.870 128.995 605.480 129.420 ;
        RECT 607.080 129.090 607.460 129.470 ;
        RECT 594.615 128.315 608.180 128.630 ;
        RECT 594.610 127.570 608.170 127.870 ;
        RECT 594.630 126.855 601.355 127.155 ;
        RECT 522.095 126.495 529.795 126.770 ;
        RECT 605.055 126.555 608.160 126.830 ;
        RECT 608.930 126.795 609.310 133.955 ;
        RECT 665.190 133.930 721.545 133.955 ;
        RECT 625.570 132.945 663.120 132.970 ;
        RECT 625.570 132.685 690.950 132.945 ;
        RECT 662.175 132.660 690.950 132.685 ;
        RECT 692.620 132.640 699.325 132.940 ;
        RECT 627.080 131.775 628.535 132.155 ;
        RECT 629.275 131.775 630.475 132.155 ;
        RECT 632.230 131.560 634.505 132.070 ;
        RECT 637.130 131.560 639.430 132.070 ;
        RECT 641.725 131.560 644.005 132.070 ;
        RECT 648.800 131.875 650.035 132.255 ;
        RECT 650.775 131.875 652.055 132.255 ;
        RECT 665.480 131.750 666.935 132.130 ;
        RECT 650.215 131.520 650.595 131.555 ;
        RECT 670.630 131.535 672.905 132.045 ;
        RECT 675.530 131.535 677.830 132.045 ;
        RECT 680.125 131.535 682.405 132.045 ;
        RECT 689.175 131.850 690.455 132.230 ;
        RECT 628.715 131.415 629.095 131.455 ;
        RECT 628.645 131.110 631.480 131.415 ;
        RECT 647.460 131.210 650.595 131.520 ;
        RECT 688.615 131.495 688.995 131.530 ;
        RECT 667.115 131.390 667.495 131.430 ;
        RECT 650.215 131.175 650.595 131.210 ;
        RECT 628.715 131.075 629.095 131.110 ;
        RECT 667.045 131.085 669.880 131.390 ;
        RECT 685.860 131.185 688.995 131.495 ;
        RECT 688.615 131.150 688.995 131.185 ;
        RECT 667.115 131.050 667.495 131.085 ;
        RECT 610.760 129.700 614.165 130.140 ;
        RECT 614.505 129.500 614.885 129.880 ;
        RECT 617.220 129.540 617.600 129.920 ;
        RECT 621.405 129.490 621.785 129.870 ;
        RECT 627.240 129.475 628.535 129.855 ;
        RECT 629.275 129.475 632.535 129.855 ;
        RECT 633.275 129.475 636.535 129.855 ;
        RECT 637.275 129.475 638.460 129.855 ;
        RECT 640.725 129.475 642.035 129.855 ;
        RECT 642.775 129.475 646.035 129.855 ;
        RECT 646.775 129.475 650.035 129.855 ;
        RECT 650.775 129.475 651.790 129.855 ;
        RECT 611.830 129.075 613.570 129.365 ;
        RECT 615.620 129.025 616.820 129.315 ;
        RECT 618.330 128.995 620.925 129.370 ;
        RECT 622.540 129.090 622.920 129.470 ;
        RECT 665.640 129.450 666.935 129.830 ;
        RECT 671.675 129.450 674.935 129.830 ;
        RECT 675.675 129.450 676.860 129.830 ;
        RECT 679.125 129.450 680.435 129.830 ;
        RECT 681.175 129.450 684.435 129.830 ;
        RECT 689.175 129.450 690.190 129.830 ;
        RECT 693.255 129.695 696.670 130.115 ;
        RECT 697.000 129.475 697.380 129.855 ;
        RECT 699.715 129.515 700.095 129.895 ;
        RECT 703.900 129.465 704.280 129.845 ;
        RECT 628.715 128.775 629.095 129.155 ;
        RECT 632.715 128.775 633.095 129.155 ;
        RECT 636.715 129.110 637.095 129.155 ;
        RECT 642.215 129.110 642.595 129.155 ;
        RECT 636.665 128.795 642.600 129.110 ;
        RECT 636.715 128.775 637.095 128.795 ;
        RECT 642.215 128.775 642.595 128.795 ;
        RECT 646.215 128.775 646.595 129.155 ;
        RECT 650.215 128.775 650.595 129.155 ;
        RECT 667.115 128.750 667.495 129.130 ;
        RECT 671.115 128.750 671.495 129.130 ;
        RECT 675.115 129.085 675.495 129.130 ;
        RECT 680.615 129.085 680.995 129.130 ;
        RECT 675.065 128.770 681.000 129.085 ;
        RECT 675.115 128.750 675.495 128.770 ;
        RECT 680.615 128.750 680.995 128.770 ;
        RECT 684.615 128.750 684.995 129.130 ;
        RECT 688.615 128.750 688.995 129.130 ;
        RECT 694.325 129.050 696.065 129.340 ;
        RECT 698.115 129.000 699.315 129.290 ;
        RECT 700.825 128.960 703.455 129.415 ;
        RECT 705.035 129.065 705.415 129.445 ;
        RECT 610.070 128.315 623.895 128.615 ;
        RECT 625.570 128.150 641.580 128.525 ;
        RECT 659.205 128.125 679.980 128.500 ;
        RECT 610.075 127.570 628.495 127.870 ;
        RECT 629.940 127.560 657.250 127.900 ;
        RECT 609.555 126.855 616.815 127.155 ;
        RECT 429.195 126.395 447.865 126.405 ;
        RECT 429.195 126.380 459.215 126.395 ;
        RECT 429.195 126.370 486.265 126.380 ;
        RECT 65.940 126.110 102.505 126.135 ;
        RECT 262.305 126.110 298.870 126.135 ;
        RECT 429.195 126.085 495.270 126.370 ;
        RECT 594.610 126.235 598.735 126.505 ;
        RECT 610.110 126.320 614.195 126.590 ;
        RECT 620.515 126.555 624.265 126.830 ;
        RECT 625.570 126.795 651.800 127.185 ;
        RECT 658.235 126.770 690.200 127.160 ;
        RECT 703.010 126.530 706.140 126.805 ;
        RECT 706.885 126.770 707.265 133.930 ;
        RECT 754.075 133.895 779.510 134.795 ;
        RECT 789.440 133.955 917.885 134.830 ;
        RECT 708.125 131.470 714.865 131.770 ;
        RECT 756.560 131.715 757.760 132.095 ;
        RECT 759.515 131.500 761.790 132.010 ;
        RECT 764.415 131.500 766.715 132.010 ;
        RECT 769.010 131.500 771.290 132.010 ;
        RECT 776.085 131.815 777.320 132.195 ;
        RECT 708.715 129.675 712.170 130.115 ;
        RECT 712.460 129.475 712.840 129.855 ;
        RECT 715.175 129.515 715.555 129.895 ;
        RECT 719.360 129.465 719.740 129.845 ;
        RECT 709.785 129.050 711.525 129.340 ;
        RECT 713.575 129.000 714.775 129.290 ;
        RECT 716.285 128.970 718.910 129.380 ;
        RECT 720.495 129.065 720.875 129.445 ;
        RECT 756.560 129.415 759.820 129.795 ;
        RECT 760.560 129.415 763.820 129.795 ;
        RECT 770.060 129.415 773.320 129.795 ;
        RECT 774.060 129.415 777.320 129.795 ;
        RECT 707.530 128.290 723.450 128.590 ;
        RECT 708.065 127.545 725.010 127.845 ;
        RECT 757.225 127.500 783.520 127.840 ;
        RECT 718.470 126.530 726.170 126.805 ;
        RECT 789.810 126.795 790.190 133.955 ;
        RECT 791.640 129.740 795.015 130.140 ;
        RECT 795.385 129.500 795.765 129.880 ;
        RECT 798.100 129.540 798.480 129.920 ;
        RECT 802.285 129.490 802.665 129.870 ;
        RECT 792.710 129.075 794.450 129.365 ;
        RECT 796.500 129.025 797.700 129.315 ;
        RECT 799.210 128.995 801.820 129.420 ;
        RECT 803.420 129.090 803.800 129.470 ;
        RECT 790.955 128.315 804.520 128.630 ;
        RECT 790.950 127.570 804.510 127.870 ;
        RECT 790.970 126.855 797.695 127.155 ;
        RECT 801.395 126.555 804.500 126.830 ;
        RECT 805.270 126.795 805.650 133.955 ;
        RECT 861.530 133.930 917.885 133.955 ;
        RECT 821.910 132.945 859.460 132.970 ;
        RECT 821.910 132.685 887.290 132.945 ;
        RECT 858.515 132.660 887.290 132.685 ;
        RECT 888.960 132.640 895.665 132.940 ;
        RECT 823.420 131.775 824.875 132.155 ;
        RECT 825.615 131.775 826.815 132.155 ;
        RECT 828.570 131.560 830.845 132.070 ;
        RECT 833.470 131.560 835.770 132.070 ;
        RECT 838.065 131.560 840.345 132.070 ;
        RECT 845.140 131.875 846.375 132.255 ;
        RECT 847.115 131.875 848.395 132.255 ;
        RECT 861.820 131.750 863.275 132.130 ;
        RECT 846.555 131.520 846.935 131.555 ;
        RECT 866.970 131.535 869.245 132.045 ;
        RECT 871.870 131.535 874.170 132.045 ;
        RECT 876.465 131.535 878.745 132.045 ;
        RECT 885.515 131.850 886.795 132.230 ;
        RECT 825.055 131.415 825.435 131.455 ;
        RECT 824.985 131.110 827.820 131.415 ;
        RECT 843.800 131.210 846.935 131.520 ;
        RECT 884.955 131.495 885.335 131.530 ;
        RECT 863.455 131.390 863.835 131.430 ;
        RECT 846.555 131.175 846.935 131.210 ;
        RECT 825.055 131.075 825.435 131.110 ;
        RECT 863.385 131.085 866.220 131.390 ;
        RECT 882.200 131.185 885.335 131.495 ;
        RECT 884.955 131.150 885.335 131.185 ;
        RECT 863.455 131.050 863.835 131.085 ;
        RECT 807.100 129.700 810.505 130.140 ;
        RECT 810.845 129.500 811.225 129.880 ;
        RECT 813.560 129.540 813.940 129.920 ;
        RECT 817.745 129.490 818.125 129.870 ;
        RECT 823.580 129.475 824.875 129.855 ;
        RECT 825.615 129.475 828.875 129.855 ;
        RECT 829.615 129.475 832.875 129.855 ;
        RECT 833.615 129.475 834.800 129.855 ;
        RECT 837.065 129.475 838.375 129.855 ;
        RECT 839.115 129.475 842.375 129.855 ;
        RECT 843.115 129.475 846.375 129.855 ;
        RECT 847.115 129.475 848.130 129.855 ;
        RECT 808.170 129.075 809.910 129.365 ;
        RECT 811.960 129.025 813.160 129.315 ;
        RECT 814.670 128.995 817.265 129.370 ;
        RECT 818.880 129.090 819.260 129.470 ;
        RECT 861.980 129.450 863.275 129.830 ;
        RECT 868.015 129.450 871.275 129.830 ;
        RECT 872.015 129.450 873.200 129.830 ;
        RECT 875.465 129.450 876.775 129.830 ;
        RECT 877.515 129.450 880.775 129.830 ;
        RECT 885.515 129.450 886.530 129.830 ;
        RECT 889.595 129.695 893.010 130.115 ;
        RECT 893.340 129.475 893.720 129.855 ;
        RECT 896.055 129.515 896.435 129.895 ;
        RECT 900.240 129.465 900.620 129.845 ;
        RECT 825.055 128.775 825.435 129.155 ;
        RECT 829.055 128.775 829.435 129.155 ;
        RECT 833.055 129.110 833.435 129.155 ;
        RECT 838.555 129.110 838.935 129.155 ;
        RECT 833.005 128.795 838.940 129.110 ;
        RECT 833.055 128.775 833.435 128.795 ;
        RECT 838.555 128.775 838.935 128.795 ;
        RECT 842.555 128.775 842.935 129.155 ;
        RECT 846.555 128.775 846.935 129.155 ;
        RECT 863.455 128.750 863.835 129.130 ;
        RECT 867.455 128.750 867.835 129.130 ;
        RECT 871.455 129.085 871.835 129.130 ;
        RECT 876.955 129.085 877.335 129.130 ;
        RECT 871.405 128.770 877.340 129.085 ;
        RECT 871.455 128.750 871.835 128.770 ;
        RECT 876.955 128.750 877.335 128.770 ;
        RECT 880.955 128.750 881.335 129.130 ;
        RECT 884.955 128.750 885.335 129.130 ;
        RECT 890.665 129.050 892.405 129.340 ;
        RECT 894.455 129.000 895.655 129.290 ;
        RECT 897.165 128.960 899.795 129.415 ;
        RECT 901.375 129.065 901.755 129.445 ;
        RECT 806.410 128.315 820.235 128.615 ;
        RECT 821.910 128.150 837.920 128.525 ;
        RECT 855.545 128.125 876.320 128.500 ;
        RECT 806.415 127.570 824.835 127.870 ;
        RECT 826.280 127.560 853.590 127.900 ;
        RECT 805.895 126.855 813.155 127.155 ;
        RECT 625.570 126.430 644.240 126.440 ;
        RECT 625.570 126.415 655.590 126.430 ;
        RECT 625.570 126.405 682.640 126.415 ;
        RECT 625.570 126.120 691.645 126.405 ;
        RECT 790.950 126.235 795.075 126.505 ;
        RECT 806.450 126.320 810.535 126.590 ;
        RECT 816.855 126.555 820.605 126.830 ;
        RECT 821.910 126.795 848.140 127.185 ;
        RECT 854.575 126.770 886.540 127.160 ;
        RECT 899.350 126.530 902.480 126.805 ;
        RECT 903.225 126.770 903.605 133.930 ;
        RECT 950.460 133.880 975.895 134.780 ;
        RECT 985.780 133.955 1114.225 134.830 ;
        RECT 904.465 131.470 911.205 131.770 ;
        RECT 952.945 131.700 954.145 132.080 ;
        RECT 955.900 131.485 958.175 131.995 ;
        RECT 960.800 131.485 963.100 131.995 ;
        RECT 965.395 131.485 967.675 131.995 ;
        RECT 972.470 131.800 973.705 132.180 ;
        RECT 905.055 129.675 908.510 130.115 ;
        RECT 908.800 129.475 909.180 129.855 ;
        RECT 911.515 129.515 911.895 129.895 ;
        RECT 915.700 129.465 916.080 129.845 ;
        RECT 906.125 129.050 907.865 129.340 ;
        RECT 909.915 129.000 911.115 129.290 ;
        RECT 912.625 128.970 915.250 129.380 ;
        RECT 916.835 129.065 917.215 129.445 ;
        RECT 952.945 129.400 956.205 129.780 ;
        RECT 956.945 129.400 960.205 129.780 ;
        RECT 966.445 129.400 969.705 129.780 ;
        RECT 970.445 129.400 973.705 129.780 ;
        RECT 903.870 128.290 919.790 128.590 ;
        RECT 904.405 127.545 921.350 127.845 ;
        RECT 953.610 127.485 979.905 127.825 ;
        RECT 914.810 126.530 922.510 126.805 ;
        RECT 986.150 126.795 986.530 133.955 ;
        RECT 987.980 129.740 991.355 130.140 ;
        RECT 991.725 129.500 992.105 129.880 ;
        RECT 994.440 129.540 994.820 129.920 ;
        RECT 998.625 129.490 999.005 129.870 ;
        RECT 989.050 129.075 990.790 129.365 ;
        RECT 992.840 129.025 994.040 129.315 ;
        RECT 995.550 128.995 998.160 129.420 ;
        RECT 999.760 129.090 1000.140 129.470 ;
        RECT 987.295 128.315 1000.860 128.630 ;
        RECT 987.290 127.570 1000.850 127.870 ;
        RECT 987.310 126.855 994.035 127.155 ;
        RECT 997.735 126.555 1000.840 126.830 ;
        RECT 1001.610 126.795 1001.990 133.955 ;
        RECT 1057.870 133.930 1114.225 133.955 ;
        RECT 1018.250 132.945 1055.800 132.970 ;
        RECT 1018.250 132.685 1083.630 132.945 ;
        RECT 1054.855 132.660 1083.630 132.685 ;
        RECT 1085.300 132.640 1092.005 132.940 ;
        RECT 1019.760 131.775 1021.215 132.155 ;
        RECT 1021.955 131.775 1023.155 132.155 ;
        RECT 1024.910 131.560 1027.185 132.070 ;
        RECT 1029.810 131.560 1032.110 132.070 ;
        RECT 1034.405 131.560 1036.685 132.070 ;
        RECT 1041.480 131.875 1042.715 132.255 ;
        RECT 1043.455 131.875 1044.735 132.255 ;
        RECT 1058.160 131.750 1059.615 132.130 ;
        RECT 1042.895 131.520 1043.275 131.555 ;
        RECT 1063.310 131.535 1065.585 132.045 ;
        RECT 1068.210 131.535 1070.510 132.045 ;
        RECT 1072.805 131.535 1075.085 132.045 ;
        RECT 1081.855 131.850 1083.135 132.230 ;
        RECT 1021.395 131.415 1021.775 131.455 ;
        RECT 1021.325 131.110 1024.160 131.415 ;
        RECT 1040.140 131.210 1043.275 131.520 ;
        RECT 1081.295 131.495 1081.675 131.530 ;
        RECT 1059.795 131.390 1060.175 131.430 ;
        RECT 1042.895 131.175 1043.275 131.210 ;
        RECT 1021.395 131.075 1021.775 131.110 ;
        RECT 1059.725 131.085 1062.560 131.390 ;
        RECT 1078.540 131.185 1081.675 131.495 ;
        RECT 1081.295 131.150 1081.675 131.185 ;
        RECT 1059.795 131.050 1060.175 131.085 ;
        RECT 1003.440 129.700 1006.845 130.140 ;
        RECT 1007.185 129.500 1007.565 129.880 ;
        RECT 1009.900 129.540 1010.280 129.920 ;
        RECT 1014.085 129.490 1014.465 129.870 ;
        RECT 1019.920 129.475 1021.215 129.855 ;
        RECT 1021.955 129.475 1025.215 129.855 ;
        RECT 1025.955 129.475 1029.215 129.855 ;
        RECT 1029.955 129.475 1031.140 129.855 ;
        RECT 1033.405 129.475 1034.715 129.855 ;
        RECT 1035.455 129.475 1038.715 129.855 ;
        RECT 1039.455 129.475 1042.715 129.855 ;
        RECT 1043.455 129.475 1044.470 129.855 ;
        RECT 1004.510 129.075 1006.250 129.365 ;
        RECT 1008.300 129.025 1009.500 129.315 ;
        RECT 1011.010 128.995 1013.605 129.370 ;
        RECT 1015.220 129.090 1015.600 129.470 ;
        RECT 1058.320 129.450 1059.615 129.830 ;
        RECT 1064.355 129.450 1067.615 129.830 ;
        RECT 1068.355 129.450 1069.540 129.830 ;
        RECT 1071.805 129.450 1073.115 129.830 ;
        RECT 1073.855 129.450 1077.115 129.830 ;
        RECT 1081.855 129.450 1082.870 129.830 ;
        RECT 1085.935 129.695 1089.350 130.115 ;
        RECT 1089.680 129.475 1090.060 129.855 ;
        RECT 1092.395 129.515 1092.775 129.895 ;
        RECT 1096.580 129.465 1096.960 129.845 ;
        RECT 1021.395 128.775 1021.775 129.155 ;
        RECT 1025.395 128.775 1025.775 129.155 ;
        RECT 1029.395 129.110 1029.775 129.155 ;
        RECT 1034.895 129.110 1035.275 129.155 ;
        RECT 1029.345 128.795 1035.280 129.110 ;
        RECT 1029.395 128.775 1029.775 128.795 ;
        RECT 1034.895 128.775 1035.275 128.795 ;
        RECT 1038.895 128.775 1039.275 129.155 ;
        RECT 1042.895 128.775 1043.275 129.155 ;
        RECT 1059.795 128.750 1060.175 129.130 ;
        RECT 1063.795 128.750 1064.175 129.130 ;
        RECT 1067.795 129.085 1068.175 129.130 ;
        RECT 1073.295 129.085 1073.675 129.130 ;
        RECT 1067.745 128.770 1073.680 129.085 ;
        RECT 1067.795 128.750 1068.175 128.770 ;
        RECT 1073.295 128.750 1073.675 128.770 ;
        RECT 1077.295 128.750 1077.675 129.130 ;
        RECT 1081.295 128.750 1081.675 129.130 ;
        RECT 1087.005 129.050 1088.745 129.340 ;
        RECT 1090.795 129.000 1091.995 129.290 ;
        RECT 1093.505 128.960 1096.135 129.415 ;
        RECT 1097.715 129.065 1098.095 129.445 ;
        RECT 1002.750 128.315 1016.575 128.615 ;
        RECT 1018.250 128.150 1034.260 128.525 ;
        RECT 1051.885 128.125 1072.660 128.500 ;
        RECT 1002.755 127.570 1021.175 127.870 ;
        RECT 1022.620 127.560 1049.930 127.900 ;
        RECT 1002.235 126.855 1009.495 127.155 ;
        RECT 821.910 126.430 840.580 126.440 ;
        RECT 821.910 126.415 851.930 126.430 ;
        RECT 821.910 126.405 878.980 126.415 ;
        RECT 821.910 126.120 887.985 126.405 ;
        RECT 987.290 126.235 991.415 126.505 ;
        RECT 1002.790 126.320 1006.875 126.590 ;
        RECT 1013.195 126.555 1016.945 126.830 ;
        RECT 1018.250 126.795 1044.480 127.185 ;
        RECT 1050.915 126.770 1082.880 127.160 ;
        RECT 1095.690 126.530 1098.820 126.805 ;
        RECT 1099.565 126.770 1099.945 133.930 ;
        RECT 1146.785 133.885 1172.220 134.785 ;
        RECT 1182.120 133.955 1310.565 134.830 ;
        RECT 1100.805 131.470 1107.545 131.770 ;
        RECT 1149.270 131.705 1150.470 132.085 ;
        RECT 1152.225 131.490 1154.500 132.000 ;
        RECT 1157.125 131.490 1159.425 132.000 ;
        RECT 1161.720 131.490 1164.000 132.000 ;
        RECT 1168.795 131.805 1170.030 132.185 ;
        RECT 1101.395 129.675 1104.850 130.115 ;
        RECT 1105.140 129.475 1105.520 129.855 ;
        RECT 1107.855 129.515 1108.235 129.895 ;
        RECT 1112.040 129.465 1112.420 129.845 ;
        RECT 1102.465 129.050 1104.205 129.340 ;
        RECT 1106.255 129.000 1107.455 129.290 ;
        RECT 1108.965 128.970 1111.590 129.380 ;
        RECT 1113.175 129.065 1113.555 129.445 ;
        RECT 1149.270 129.405 1152.530 129.785 ;
        RECT 1153.270 129.405 1156.530 129.785 ;
        RECT 1162.770 129.405 1166.030 129.785 ;
        RECT 1166.770 129.405 1170.030 129.785 ;
        RECT 1100.210 128.290 1116.130 128.590 ;
        RECT 1100.745 127.545 1117.690 127.845 ;
        RECT 1149.935 127.490 1176.230 127.830 ;
        RECT 1111.150 126.530 1118.850 126.805 ;
        RECT 1182.490 126.795 1182.870 133.955 ;
        RECT 1184.320 129.740 1187.695 130.140 ;
        RECT 1188.065 129.500 1188.445 129.880 ;
        RECT 1190.780 129.540 1191.160 129.920 ;
        RECT 1194.965 129.490 1195.345 129.870 ;
        RECT 1185.390 129.075 1187.130 129.365 ;
        RECT 1189.180 129.025 1190.380 129.315 ;
        RECT 1191.890 128.995 1194.500 129.420 ;
        RECT 1196.100 129.090 1196.480 129.470 ;
        RECT 1183.635 128.315 1197.200 128.630 ;
        RECT 1183.630 127.570 1197.190 127.870 ;
        RECT 1183.650 126.855 1190.375 127.155 ;
        RECT 1194.075 126.555 1197.180 126.830 ;
        RECT 1197.950 126.795 1198.330 133.955 ;
        RECT 1254.210 133.930 1310.565 133.955 ;
        RECT 1214.590 132.945 1252.140 132.970 ;
        RECT 1214.590 132.685 1279.970 132.945 ;
        RECT 1251.195 132.660 1279.970 132.685 ;
        RECT 1281.640 132.640 1288.345 132.940 ;
        RECT 1216.100 131.775 1217.555 132.155 ;
        RECT 1218.295 131.775 1219.495 132.155 ;
        RECT 1221.250 131.560 1223.525 132.070 ;
        RECT 1226.150 131.560 1228.450 132.070 ;
        RECT 1230.745 131.560 1233.025 132.070 ;
        RECT 1237.820 131.875 1239.055 132.255 ;
        RECT 1239.795 131.875 1241.075 132.255 ;
        RECT 1254.500 131.750 1255.955 132.130 ;
        RECT 1256.695 131.750 1257.895 132.130 ;
        RECT 1239.235 131.520 1239.615 131.555 ;
        RECT 1259.650 131.535 1261.925 132.045 ;
        RECT 1264.550 131.535 1266.850 132.045 ;
        RECT 1269.145 131.535 1271.425 132.045 ;
        RECT 1276.220 131.850 1277.455 132.230 ;
        RECT 1278.195 131.850 1279.475 132.230 ;
        RECT 1217.735 131.415 1218.115 131.455 ;
        RECT 1217.665 131.110 1220.500 131.415 ;
        RECT 1236.480 131.210 1239.615 131.520 ;
        RECT 1277.635 131.495 1278.015 131.530 ;
        RECT 1256.135 131.390 1256.515 131.430 ;
        RECT 1239.235 131.175 1239.615 131.210 ;
        RECT 1217.735 131.075 1218.115 131.110 ;
        RECT 1256.065 131.085 1258.900 131.390 ;
        RECT 1274.880 131.185 1278.015 131.495 ;
        RECT 1277.635 131.150 1278.015 131.185 ;
        RECT 1256.135 131.050 1256.515 131.085 ;
        RECT 1199.780 129.700 1203.185 130.140 ;
        RECT 1203.525 129.500 1203.905 129.880 ;
        RECT 1206.240 129.540 1206.620 129.920 ;
        RECT 1210.425 129.490 1210.805 129.870 ;
        RECT 1216.260 129.475 1217.555 129.855 ;
        RECT 1218.295 129.475 1221.555 129.855 ;
        RECT 1222.295 129.475 1225.555 129.855 ;
        RECT 1226.295 129.475 1227.480 129.855 ;
        RECT 1229.745 129.475 1231.055 129.855 ;
        RECT 1231.795 129.475 1235.055 129.855 ;
        RECT 1235.795 129.475 1239.055 129.855 ;
        RECT 1239.795 129.475 1240.810 129.855 ;
        RECT 1200.850 129.075 1202.590 129.365 ;
        RECT 1204.640 129.025 1205.840 129.315 ;
        RECT 1207.350 128.995 1209.945 129.370 ;
        RECT 1211.560 129.090 1211.940 129.470 ;
        RECT 1254.660 129.450 1255.955 129.830 ;
        RECT 1256.695 129.450 1259.955 129.830 ;
        RECT 1260.695 129.450 1263.955 129.830 ;
        RECT 1264.695 129.450 1265.880 129.830 ;
        RECT 1268.145 129.450 1269.455 129.830 ;
        RECT 1270.195 129.450 1273.455 129.830 ;
        RECT 1274.195 129.450 1277.455 129.830 ;
        RECT 1278.195 129.450 1279.210 129.830 ;
        RECT 1282.275 129.695 1285.690 130.115 ;
        RECT 1286.020 129.475 1286.400 129.855 ;
        RECT 1288.735 129.515 1289.115 129.895 ;
        RECT 1292.920 129.465 1293.300 129.845 ;
        RECT 1217.735 128.775 1218.115 129.155 ;
        RECT 1221.735 128.775 1222.115 129.155 ;
        RECT 1225.735 129.110 1226.115 129.155 ;
        RECT 1231.235 129.110 1231.615 129.155 ;
        RECT 1225.685 128.795 1231.620 129.110 ;
        RECT 1225.735 128.775 1226.115 128.795 ;
        RECT 1231.235 128.775 1231.615 128.795 ;
        RECT 1235.235 128.775 1235.615 129.155 ;
        RECT 1239.235 128.775 1239.615 129.155 ;
        RECT 1256.135 128.750 1256.515 129.130 ;
        RECT 1260.135 128.750 1260.515 129.130 ;
        RECT 1264.135 129.085 1264.515 129.130 ;
        RECT 1269.635 129.085 1270.015 129.130 ;
        RECT 1264.085 128.770 1270.020 129.085 ;
        RECT 1264.135 128.750 1264.515 128.770 ;
        RECT 1269.635 128.750 1270.015 128.770 ;
        RECT 1273.635 128.750 1274.015 129.130 ;
        RECT 1277.635 128.750 1278.015 129.130 ;
        RECT 1283.345 129.050 1285.085 129.340 ;
        RECT 1287.135 129.000 1288.335 129.290 ;
        RECT 1289.845 128.960 1292.475 129.415 ;
        RECT 1294.055 129.065 1294.435 129.445 ;
        RECT 1199.090 128.315 1212.915 128.615 ;
        RECT 1214.590 128.150 1230.600 128.525 ;
        RECT 1248.225 128.125 1269.000 128.500 ;
        RECT 1281.625 128.290 1295.240 128.590 ;
        RECT 1199.095 127.570 1217.515 127.870 ;
        RECT 1218.960 127.560 1246.270 127.900 ;
        RECT 1257.360 127.535 1279.915 127.875 ;
        RECT 1281.025 127.545 1295.670 127.845 ;
        RECT 1198.575 126.855 1205.835 127.155 ;
        RECT 1018.250 126.430 1036.920 126.440 ;
        RECT 1018.250 126.415 1048.270 126.430 ;
        RECT 1018.250 126.405 1075.320 126.415 ;
        RECT 1018.250 126.120 1084.325 126.405 ;
        RECT 1183.630 126.235 1187.755 126.505 ;
        RECT 1199.130 126.320 1203.215 126.590 ;
        RECT 1209.535 126.555 1213.285 126.830 ;
        RECT 1214.590 126.795 1240.820 127.185 ;
        RECT 1247.255 126.770 1279.220 127.160 ;
        RECT 1292.030 126.530 1295.160 126.805 ;
        RECT 1295.905 126.770 1296.285 133.930 ;
        RECT 1297.145 131.470 1303.885 131.770 ;
        RECT 1297.735 129.675 1301.190 130.115 ;
        RECT 1304.195 129.515 1304.575 129.895 ;
        RECT 1302.595 129.000 1303.795 129.290 ;
        RECT 1309.515 129.065 1309.895 129.445 ;
        RECT 1296.550 128.290 1312.470 128.590 ;
        RECT 1297.085 127.545 1314.030 127.845 ;
        RECT 1214.590 126.430 1233.260 126.440 ;
        RECT 1214.590 126.415 1244.610 126.430 ;
        RECT 1214.590 126.405 1271.660 126.415 ;
        RECT 1214.590 126.120 1280.665 126.405 ;
        RECT 655.080 126.095 691.645 126.120 ;
        RECT 851.420 126.095 887.985 126.120 ;
        RECT 1047.760 126.095 1084.325 126.120 ;
        RECT 1244.100 126.095 1280.665 126.120 ;
        RECT 458.705 126.060 495.270 126.085 ;
        RECT 6.705 125.675 10.835 125.975 ;
        RECT -59.625 124.780 -56.060 124.790 ;
        RECT -59.625 124.455 -55.265 124.780 ;
        RECT -9.300 124.535 -3.385 124.870 ;
        RECT -6.030 124.515 -3.385 124.535 ;
        RECT -56.220 124.445 -55.265 124.455 ;
        RECT -79.030 123.815 -75.730 124.195 ;
        RECT -75.030 123.815 -71.730 124.195 ;
        RECT -65.530 123.815 -62.230 124.195 ;
        RECT -61.530 123.815 -58.230 124.195 ;
        RECT -28.705 123.895 -25.405 124.275 ;
        RECT -24.705 123.895 -21.405 124.275 ;
        RECT -15.205 123.895 -11.905 124.275 ;
        RECT -11.205 123.895 -7.905 124.275 ;
        RECT -79.030 121.815 -77.745 122.195 ;
        RECT -59.715 121.815 -58.230 122.195 ;
        RECT -28.705 121.895 -27.420 122.275 ;
        RECT -9.390 121.895 -7.905 122.275 ;
        RECT -77.525 121.135 -76.005 121.495 ;
        RECT -27.200 121.215 -25.680 121.575 ;
        RECT 4.330 119.845 4.710 125.675 ;
        RECT 13.210 125.625 17.710 125.935 ;
        RECT 22.165 125.675 26.295 125.975 ;
        RECT 9.170 125.075 15.560 125.365 ;
        RECT 8.585 124.495 19.240 124.830 ;
        RECT 7.935 123.910 10.855 124.210 ;
        RECT 14.400 123.895 17.770 124.195 ;
        RECT 6.150 123.160 6.530 123.540 ;
        RECT 8.555 123.175 10.335 123.465 ;
        RECT 11.810 123.265 13.000 123.550 ;
        RECT 15.930 123.145 17.240 123.465 ;
        RECT 7.285 122.560 7.665 122.940 ;
        RECT 11.030 122.600 11.410 122.980 ;
        RECT 13.740 122.590 14.120 122.970 ;
        RECT 15.150 122.435 18.330 122.755 ;
        RECT 5.080 119.845 9.175 119.850 ;
        RECT 19.790 119.845 20.170 125.675 ;
        RECT 28.670 125.625 33.170 125.935 ;
        RECT 120.120 125.650 124.250 125.950 ;
        RECT 35.900 125.440 71.810 125.465 ;
        RECT 24.630 125.075 31.020 125.365 ;
        RECT 35.900 125.195 102.905 125.440 ;
        RECT 71.160 125.170 102.905 125.195 ;
        RECT 107.125 125.050 113.515 125.340 ;
        RECT 24.045 124.495 34.550 124.830 ;
        RECT 59.520 124.630 70.070 124.965 ;
        RECT 106.540 124.470 117.020 124.805 ;
        RECT 23.395 123.910 26.315 124.210 ;
        RECT 29.860 123.895 33.230 124.195 ;
        RECT 38.110 123.990 39.415 124.370 ;
        RECT 40.115 123.990 43.415 124.370 ;
        RECT 44.115 123.990 47.415 124.370 ;
        RECT 48.115 123.990 49.475 124.370 ;
        RECT 51.450 123.990 52.915 124.370 ;
        RECT 53.615 123.990 56.915 124.370 ;
        RECT 57.615 123.990 60.915 124.370 ;
        RECT 61.615 123.990 62.795 124.370 ;
        RECT 76.510 123.965 77.815 124.345 ;
        RECT 82.515 123.965 85.815 124.345 ;
        RECT 86.515 123.965 87.875 124.345 ;
        RECT 89.850 123.965 91.315 124.345 ;
        RECT 92.015 123.965 95.315 124.345 ;
        RECT 100.015 123.965 101.195 124.345 ;
        RECT 39.575 123.645 39.955 123.680 ;
        RECT 21.610 123.160 21.990 123.540 ;
        RECT 24.015 123.175 25.795 123.465 ;
        RECT 27.270 123.265 28.460 123.550 ;
        RECT 31.390 123.145 32.700 123.465 ;
        RECT 39.310 123.335 42.320 123.645 ;
        RECT 39.575 123.300 39.955 123.335 ;
        RECT 43.575 123.300 44.665 123.680 ;
        RECT 47.575 123.675 47.955 123.680 ;
        RECT 45.095 123.310 47.960 123.675 ;
        RECT 53.075 123.655 53.455 123.680 ;
        RECT 53.060 123.335 55.205 123.655 ;
        RECT 47.575 123.300 47.955 123.310 ;
        RECT 53.075 123.300 53.455 123.335 ;
        RECT 56.120 123.300 57.455 123.680 ;
        RECT 61.075 123.660 61.455 123.680 ;
        RECT 58.610 123.340 61.520 123.660 ;
        RECT 77.975 123.620 78.355 123.655 ;
        RECT 61.075 123.300 61.455 123.340 ;
        RECT 77.710 123.310 80.720 123.620 ;
        RECT 77.975 123.275 78.355 123.310 ;
        RECT 81.975 123.275 83.065 123.655 ;
        RECT 85.975 123.650 86.355 123.655 ;
        RECT 83.495 123.285 86.360 123.650 ;
        RECT 91.475 123.630 91.855 123.655 ;
        RECT 91.460 123.310 93.605 123.630 ;
        RECT 85.975 123.275 86.355 123.285 ;
        RECT 91.475 123.275 91.855 123.310 ;
        RECT 94.520 123.275 95.855 123.655 ;
        RECT 99.475 123.635 99.855 123.655 ;
        RECT 97.010 123.315 99.920 123.635 ;
        RECT 99.475 123.275 99.855 123.315 ;
        RECT 104.105 123.135 104.485 123.515 ;
        RECT 106.510 123.150 108.290 123.440 ;
        RECT 109.765 123.240 110.955 123.525 ;
        RECT 113.885 123.120 115.195 123.440 ;
        RECT 22.745 122.560 23.125 122.940 ;
        RECT 26.490 122.600 26.870 122.980 ;
        RECT 29.200 122.590 29.580 122.970 ;
        RECT 30.610 122.435 33.790 122.755 ;
        RECT 105.240 122.535 105.620 122.915 ;
        RECT 108.985 122.575 109.365 122.955 ;
        RECT 111.695 122.565 112.075 122.945 ;
        RECT 113.105 122.410 116.285 122.730 ;
        RECT 37.925 121.990 39.415 122.370 ;
        RECT 40.115 121.990 41.400 122.370 ;
        RECT 59.430 121.990 60.915 122.370 ;
        RECT 61.615 121.990 62.690 122.370 ;
        RECT 76.325 121.965 77.815 122.345 ;
        RECT 100.015 121.965 101.090 122.345 ;
        RECT 39.575 121.300 40.665 121.680 ;
        RECT 41.620 121.310 43.140 121.670 ;
        RECT 44.060 121.305 56.910 121.640 ;
        RECT 61.075 121.635 61.455 121.680 ;
        RECT 60.340 121.335 61.650 121.635 ;
        RECT 61.075 121.300 61.455 121.335 ;
        RECT 77.975 121.275 79.065 121.655 ;
        RECT 80.020 121.285 81.540 121.645 ;
        RECT 82.460 121.280 95.310 121.615 ;
        RECT 99.475 121.610 99.855 121.655 ;
        RECT 98.740 121.310 100.050 121.610 ;
        RECT 99.475 121.275 99.855 121.310 ;
        RECT 36.430 120.780 69.510 120.790 ;
        RECT 36.430 120.440 101.485 120.780 ;
        RECT 68.535 120.415 101.485 120.440 ;
        RECT 103.280 120.405 107.540 120.760 ;
        RECT 20.540 119.845 24.635 119.850 ;
        RECT 3.960 119.840 9.175 119.845 ;
        RECT 19.420 119.840 24.635 119.845 ;
        RECT 34.880 119.840 75.130 119.845 ;
        RECT 3.960 119.820 75.130 119.840 ;
        RECT 101.485 119.820 107.130 119.825 ;
        RECT 117.745 119.820 118.125 125.650 ;
        RECT 126.625 125.600 131.125 125.910 ;
        RECT 203.070 125.675 207.200 125.975 ;
        RECT 122.585 125.050 128.975 125.340 ;
        RECT 122.000 124.470 138.020 124.805 ;
        RECT 186.870 124.545 192.785 124.880 ;
        RECT 190.140 124.525 192.785 124.545 ;
        RECT 121.350 123.885 124.270 124.185 ;
        RECT 127.815 123.870 131.185 124.170 ;
        RECT 167.465 123.905 170.765 124.285 ;
        RECT 171.465 123.905 174.765 124.285 ;
        RECT 180.965 123.905 184.265 124.285 ;
        RECT 184.965 123.905 188.265 124.285 ;
        RECT 119.565 123.135 119.945 123.515 ;
        RECT 121.970 123.150 123.750 123.440 ;
        RECT 125.225 123.240 126.415 123.525 ;
        RECT 129.345 123.120 130.655 123.440 ;
        RECT 120.700 122.535 121.080 122.915 ;
        RECT 124.445 122.575 124.825 122.955 ;
        RECT 127.155 122.565 127.535 122.945 ;
        RECT 128.565 122.410 131.745 122.730 ;
        RECT 167.465 121.905 168.750 122.285 ;
        RECT 186.780 121.905 188.265 122.285 ;
        RECT 118.845 121.325 122.995 121.595 ;
        RECT 168.970 121.225 170.490 121.585 ;
        RECT 200.695 119.845 201.075 125.675 ;
        RECT 209.575 125.625 214.075 125.935 ;
        RECT 218.530 125.675 222.660 125.975 ;
        RECT 205.535 125.075 211.925 125.365 ;
        RECT 204.950 124.495 215.605 124.830 ;
        RECT 204.300 123.910 207.220 124.210 ;
        RECT 210.765 123.895 214.135 124.195 ;
        RECT 202.515 123.160 202.895 123.540 ;
        RECT 204.920 123.175 206.700 123.465 ;
        RECT 208.175 123.265 209.365 123.550 ;
        RECT 212.295 123.145 213.605 123.465 ;
        RECT 203.650 122.560 204.030 122.940 ;
        RECT 207.395 122.600 207.775 122.980 ;
        RECT 210.105 122.590 210.485 122.970 ;
        RECT 211.515 122.435 214.695 122.755 ;
        RECT 201.445 119.845 205.540 119.850 ;
        RECT 216.155 119.845 216.535 125.675 ;
        RECT 225.035 125.625 229.535 125.935 ;
        RECT 316.485 125.650 320.615 125.950 ;
        RECT 232.265 125.440 268.175 125.465 ;
        RECT 220.995 125.075 227.385 125.365 ;
        RECT 232.265 125.195 299.270 125.440 ;
        RECT 267.525 125.170 299.270 125.195 ;
        RECT 303.490 125.050 309.880 125.340 ;
        RECT 220.410 124.495 230.915 124.830 ;
        RECT 255.885 124.630 266.435 124.965 ;
        RECT 302.905 124.470 313.385 124.805 ;
        RECT 219.760 123.910 222.680 124.210 ;
        RECT 226.225 123.895 229.595 124.195 ;
        RECT 234.475 123.990 235.780 124.370 ;
        RECT 236.480 123.990 239.780 124.370 ;
        RECT 240.480 123.990 243.780 124.370 ;
        RECT 244.480 123.990 245.840 124.370 ;
        RECT 247.815 123.990 249.280 124.370 ;
        RECT 249.980 123.990 253.280 124.370 ;
        RECT 253.980 123.990 257.280 124.370 ;
        RECT 257.980 123.990 259.160 124.370 ;
        RECT 272.875 123.965 274.180 124.345 ;
        RECT 278.880 123.965 282.180 124.345 ;
        RECT 282.880 123.965 284.240 124.345 ;
        RECT 286.215 123.965 287.680 124.345 ;
        RECT 288.380 123.965 291.680 124.345 ;
        RECT 296.380 123.965 297.560 124.345 ;
        RECT 235.940 123.645 236.320 123.680 ;
        RECT 217.975 123.160 218.355 123.540 ;
        RECT 220.380 123.175 222.160 123.465 ;
        RECT 223.635 123.265 224.825 123.550 ;
        RECT 227.755 123.145 229.065 123.465 ;
        RECT 235.675 123.335 238.685 123.645 ;
        RECT 235.940 123.300 236.320 123.335 ;
        RECT 239.940 123.300 241.030 123.680 ;
        RECT 243.940 123.675 244.320 123.680 ;
        RECT 241.460 123.310 244.325 123.675 ;
        RECT 249.440 123.655 249.820 123.680 ;
        RECT 249.425 123.335 251.570 123.655 ;
        RECT 243.940 123.300 244.320 123.310 ;
        RECT 249.440 123.300 249.820 123.335 ;
        RECT 252.485 123.300 253.820 123.680 ;
        RECT 257.440 123.660 257.820 123.680 ;
        RECT 254.975 123.340 257.885 123.660 ;
        RECT 274.340 123.620 274.720 123.655 ;
        RECT 257.440 123.300 257.820 123.340 ;
        RECT 274.075 123.310 277.085 123.620 ;
        RECT 274.340 123.275 274.720 123.310 ;
        RECT 278.340 123.275 279.430 123.655 ;
        RECT 282.340 123.650 282.720 123.655 ;
        RECT 279.860 123.285 282.725 123.650 ;
        RECT 287.840 123.630 288.220 123.655 ;
        RECT 287.825 123.310 289.970 123.630 ;
        RECT 282.340 123.275 282.720 123.285 ;
        RECT 287.840 123.275 288.220 123.310 ;
        RECT 290.885 123.275 292.220 123.655 ;
        RECT 295.840 123.635 296.220 123.655 ;
        RECT 293.375 123.315 296.285 123.635 ;
        RECT 295.840 123.275 296.220 123.315 ;
        RECT 300.470 123.135 300.850 123.515 ;
        RECT 302.875 123.150 304.655 123.440 ;
        RECT 306.130 123.240 307.320 123.525 ;
        RECT 310.250 123.120 311.560 123.440 ;
        RECT 219.110 122.560 219.490 122.940 ;
        RECT 222.855 122.600 223.235 122.980 ;
        RECT 225.565 122.590 225.945 122.970 ;
        RECT 226.975 122.435 230.155 122.755 ;
        RECT 301.605 122.535 301.985 122.915 ;
        RECT 305.350 122.575 305.730 122.955 ;
        RECT 308.060 122.565 308.440 122.945 ;
        RECT 309.470 122.410 312.650 122.730 ;
        RECT 234.290 121.990 235.780 122.370 ;
        RECT 236.480 121.990 237.765 122.370 ;
        RECT 255.795 121.990 257.280 122.370 ;
        RECT 257.980 121.990 259.055 122.370 ;
        RECT 272.690 121.965 274.180 122.345 ;
        RECT 296.380 121.965 297.455 122.345 ;
        RECT 235.940 121.300 237.030 121.680 ;
        RECT 237.985 121.310 239.505 121.670 ;
        RECT 240.425 121.305 253.275 121.640 ;
        RECT 257.440 121.635 257.820 121.680 ;
        RECT 256.705 121.335 258.015 121.635 ;
        RECT 257.440 121.300 257.820 121.335 ;
        RECT 274.340 121.275 275.430 121.655 ;
        RECT 276.385 121.285 277.905 121.645 ;
        RECT 278.825 121.280 291.675 121.615 ;
        RECT 295.840 121.610 296.220 121.655 ;
        RECT 295.105 121.310 296.415 121.610 ;
        RECT 295.840 121.275 296.220 121.310 ;
        RECT 232.795 120.780 265.875 120.790 ;
        RECT 232.795 120.440 297.850 120.780 ;
        RECT 264.900 120.415 297.850 120.440 ;
        RECT 299.645 120.405 303.905 120.760 ;
        RECT 216.905 119.845 221.000 119.850 ;
        RECT 200.325 119.840 205.540 119.845 ;
        RECT 215.785 119.840 221.000 119.845 ;
        RECT 231.245 119.840 271.495 119.845 ;
        RECT 118.495 119.820 122.590 119.825 ;
        RECT 3.960 119.815 107.130 119.820 ;
        RECT 117.375 119.815 122.590 119.820 ;
        RECT 200.325 119.820 271.495 119.840 ;
        RECT 297.850 119.820 303.495 119.825 ;
        RECT 314.110 119.820 314.490 125.650 ;
        RECT 322.990 125.600 327.490 125.910 ;
        RECT 399.470 125.625 403.600 125.925 ;
        RECT 318.950 125.050 325.340 125.340 ;
        RECT 318.365 124.470 334.385 124.805 ;
        RECT 383.260 124.505 389.175 124.840 ;
        RECT 386.530 124.485 389.175 124.505 ;
        RECT 317.715 123.885 320.635 124.185 ;
        RECT 324.180 123.870 327.550 124.170 ;
        RECT 363.855 123.865 367.155 124.245 ;
        RECT 367.855 123.865 371.155 124.245 ;
        RECT 377.355 123.865 380.655 124.245 ;
        RECT 381.355 123.865 384.655 124.245 ;
        RECT 315.930 123.135 316.310 123.515 ;
        RECT 318.335 123.150 320.115 123.440 ;
        RECT 321.590 123.240 322.780 123.525 ;
        RECT 325.710 123.120 327.020 123.440 ;
        RECT 317.065 122.535 317.445 122.915 ;
        RECT 320.810 122.575 321.190 122.955 ;
        RECT 323.520 122.565 323.900 122.945 ;
        RECT 324.930 122.410 328.110 122.730 ;
        RECT 363.855 121.865 365.140 122.245 ;
        RECT 383.170 121.865 384.655 122.245 ;
        RECT 315.210 121.325 319.360 121.595 ;
        RECT 365.360 121.185 366.880 121.545 ;
        RECT 314.860 119.820 318.955 119.825 ;
        RECT 200.325 119.815 303.495 119.820 ;
        RECT 313.740 119.815 318.955 119.820 ;
        RECT -82.715 118.770 -56.060 119.670 ;
        RECT -32.390 118.850 -5.735 119.750 ;
        RECT 3.960 118.945 132.405 119.815 ;
        RECT 74.830 118.920 132.405 118.945 ;
        RECT 163.780 118.860 190.435 119.760 ;
        RECT 200.325 118.945 328.770 119.815 ;
        RECT 397.095 119.795 397.475 125.625 ;
        RECT 405.975 125.575 410.475 125.885 ;
        RECT 414.930 125.625 419.060 125.925 ;
        RECT 401.935 125.025 408.325 125.315 ;
        RECT 401.350 124.445 412.005 124.780 ;
        RECT 400.700 123.860 403.620 124.160 ;
        RECT 407.165 123.845 410.535 124.145 ;
        RECT 398.915 123.110 399.295 123.490 ;
        RECT 401.320 123.125 403.100 123.415 ;
        RECT 404.575 123.215 405.765 123.500 ;
        RECT 408.695 123.095 410.005 123.415 ;
        RECT 400.050 122.510 400.430 122.890 ;
        RECT 403.795 122.550 404.175 122.930 ;
        RECT 406.505 122.540 406.885 122.920 ;
        RECT 407.915 122.385 411.095 122.705 ;
        RECT 397.845 119.795 401.940 119.800 ;
        RECT 412.555 119.795 412.935 125.625 ;
        RECT 421.435 125.575 425.935 125.885 ;
        RECT 512.885 125.600 517.015 125.900 ;
        RECT 428.665 125.390 464.575 125.415 ;
        RECT 417.395 125.025 423.785 125.315 ;
        RECT 428.665 125.145 495.670 125.390 ;
        RECT 463.925 125.120 495.670 125.145 ;
        RECT 499.890 125.000 506.280 125.290 ;
        RECT 416.810 124.445 427.315 124.780 ;
        RECT 452.285 124.580 462.835 124.915 ;
        RECT 499.305 124.420 509.785 124.755 ;
        RECT 416.160 123.860 419.080 124.160 ;
        RECT 422.625 123.845 425.995 124.145 ;
        RECT 430.875 123.940 432.180 124.320 ;
        RECT 432.880 123.940 436.180 124.320 ;
        RECT 436.880 123.940 440.180 124.320 ;
        RECT 440.880 123.940 442.240 124.320 ;
        RECT 444.215 123.940 445.680 124.320 ;
        RECT 446.380 123.940 449.680 124.320 ;
        RECT 450.380 123.940 453.680 124.320 ;
        RECT 454.380 123.940 455.560 124.320 ;
        RECT 469.275 123.915 470.580 124.295 ;
        RECT 475.280 123.915 478.580 124.295 ;
        RECT 479.280 123.915 480.640 124.295 ;
        RECT 482.615 123.915 484.080 124.295 ;
        RECT 484.780 123.915 488.080 124.295 ;
        RECT 492.780 123.915 493.960 124.295 ;
        RECT 432.340 123.595 432.720 123.630 ;
        RECT 414.375 123.110 414.755 123.490 ;
        RECT 416.780 123.125 418.560 123.415 ;
        RECT 420.035 123.215 421.225 123.500 ;
        RECT 424.155 123.095 425.465 123.415 ;
        RECT 432.075 123.285 435.085 123.595 ;
        RECT 432.340 123.250 432.720 123.285 ;
        RECT 436.340 123.250 437.430 123.630 ;
        RECT 440.340 123.625 440.720 123.630 ;
        RECT 437.860 123.260 440.725 123.625 ;
        RECT 445.840 123.605 446.220 123.630 ;
        RECT 445.825 123.285 447.970 123.605 ;
        RECT 440.340 123.250 440.720 123.260 ;
        RECT 445.840 123.250 446.220 123.285 ;
        RECT 448.885 123.250 450.220 123.630 ;
        RECT 453.840 123.610 454.220 123.630 ;
        RECT 451.375 123.290 454.285 123.610 ;
        RECT 470.740 123.570 471.120 123.605 ;
        RECT 453.840 123.250 454.220 123.290 ;
        RECT 470.475 123.260 473.485 123.570 ;
        RECT 470.740 123.225 471.120 123.260 ;
        RECT 474.740 123.225 475.830 123.605 ;
        RECT 478.740 123.600 479.120 123.605 ;
        RECT 476.260 123.235 479.125 123.600 ;
        RECT 484.240 123.580 484.620 123.605 ;
        RECT 484.225 123.260 486.370 123.580 ;
        RECT 478.740 123.225 479.120 123.235 ;
        RECT 484.240 123.225 484.620 123.260 ;
        RECT 487.285 123.225 488.620 123.605 ;
        RECT 492.240 123.585 492.620 123.605 ;
        RECT 489.775 123.265 492.685 123.585 ;
        RECT 492.240 123.225 492.620 123.265 ;
        RECT 496.870 123.085 497.250 123.465 ;
        RECT 499.275 123.100 501.055 123.390 ;
        RECT 502.530 123.190 503.720 123.475 ;
        RECT 506.650 123.070 507.960 123.390 ;
        RECT 415.510 122.510 415.890 122.890 ;
        RECT 419.255 122.550 419.635 122.930 ;
        RECT 421.965 122.540 422.345 122.920 ;
        RECT 423.375 122.385 426.555 122.705 ;
        RECT 498.005 122.485 498.385 122.865 ;
        RECT 501.750 122.525 502.130 122.905 ;
        RECT 504.460 122.515 504.840 122.895 ;
        RECT 505.870 122.360 509.050 122.680 ;
        RECT 430.690 121.940 432.180 122.320 ;
        RECT 432.880 121.940 434.165 122.320 ;
        RECT 452.195 121.940 453.680 122.320 ;
        RECT 454.380 121.940 455.455 122.320 ;
        RECT 469.090 121.915 470.580 122.295 ;
        RECT 492.780 121.915 493.855 122.295 ;
        RECT 432.340 121.250 433.430 121.630 ;
        RECT 434.385 121.260 435.905 121.620 ;
        RECT 436.825 121.255 449.675 121.590 ;
        RECT 453.840 121.585 454.220 121.630 ;
        RECT 453.105 121.285 454.415 121.585 ;
        RECT 453.840 121.250 454.220 121.285 ;
        RECT 470.740 121.225 471.830 121.605 ;
        RECT 472.785 121.235 474.305 121.595 ;
        RECT 475.225 121.230 488.075 121.565 ;
        RECT 492.240 121.560 492.620 121.605 ;
        RECT 491.505 121.260 492.815 121.560 ;
        RECT 492.240 121.225 492.620 121.260 ;
        RECT 429.195 120.730 462.275 120.740 ;
        RECT 429.195 120.390 494.250 120.730 ;
        RECT 461.300 120.365 494.250 120.390 ;
        RECT 496.045 120.355 500.305 120.710 ;
        RECT 413.305 119.795 417.400 119.800 ;
        RECT 396.725 119.790 401.940 119.795 ;
        RECT 412.185 119.790 417.400 119.795 ;
        RECT 427.645 119.790 467.895 119.795 ;
        RECT 396.725 119.770 467.895 119.790 ;
        RECT 494.250 119.770 499.895 119.775 ;
        RECT 510.510 119.770 510.890 125.600 ;
        RECT 519.390 125.550 523.890 125.860 ;
        RECT 595.845 125.660 599.975 125.960 ;
        RECT 515.350 125.000 521.740 125.290 ;
        RECT 514.765 124.420 530.785 124.755 ;
        RECT 579.580 124.550 585.495 124.885 ;
        RECT 582.850 124.530 585.495 124.550 ;
        RECT 514.115 123.835 517.035 124.135 ;
        RECT 520.580 123.820 523.950 124.120 ;
        RECT 560.175 123.910 563.475 124.290 ;
        RECT 564.175 123.910 567.475 124.290 ;
        RECT 573.675 123.910 576.975 124.290 ;
        RECT 577.675 123.910 580.975 124.290 ;
        RECT 512.330 123.085 512.710 123.465 ;
        RECT 514.735 123.100 516.515 123.390 ;
        RECT 517.990 123.190 519.180 123.475 ;
        RECT 522.110 123.070 523.420 123.390 ;
        RECT 513.465 122.485 513.845 122.865 ;
        RECT 517.210 122.525 517.590 122.905 ;
        RECT 519.920 122.515 520.300 122.895 ;
        RECT 521.330 122.360 524.510 122.680 ;
        RECT 560.175 121.910 561.460 122.290 ;
        RECT 579.490 121.910 580.975 122.290 ;
        RECT 511.610 121.275 515.760 121.545 ;
        RECT 561.680 121.230 563.200 121.590 ;
        RECT 593.470 119.830 593.850 125.660 ;
        RECT 602.350 125.610 606.850 125.920 ;
        RECT 611.305 125.660 615.435 125.960 ;
        RECT 598.310 125.060 604.700 125.350 ;
        RECT 597.725 124.480 608.380 124.815 ;
        RECT 597.075 123.895 599.995 124.195 ;
        RECT 603.540 123.880 606.910 124.180 ;
        RECT 595.290 123.145 595.670 123.525 ;
        RECT 597.695 123.160 599.475 123.450 ;
        RECT 600.950 123.250 602.140 123.535 ;
        RECT 605.070 123.130 606.380 123.450 ;
        RECT 596.425 122.545 596.805 122.925 ;
        RECT 600.170 122.585 600.550 122.965 ;
        RECT 602.880 122.575 603.260 122.955 ;
        RECT 604.290 122.420 607.470 122.740 ;
        RECT 594.220 119.830 598.315 119.835 ;
        RECT 608.930 119.830 609.310 125.660 ;
        RECT 617.810 125.610 622.310 125.920 ;
        RECT 709.260 125.635 713.390 125.935 ;
        RECT 625.040 125.425 660.950 125.450 ;
        RECT 613.770 125.060 620.160 125.350 ;
        RECT 625.040 125.180 692.045 125.425 ;
        RECT 660.300 125.155 692.045 125.180 ;
        RECT 696.265 125.035 702.655 125.325 ;
        RECT 613.185 124.480 623.690 124.815 ;
        RECT 648.660 124.615 659.210 124.950 ;
        RECT 695.680 124.455 706.160 124.790 ;
        RECT 612.535 123.895 615.455 124.195 ;
        RECT 619.000 123.880 622.370 124.180 ;
        RECT 627.250 123.975 628.555 124.355 ;
        RECT 629.255 123.975 632.555 124.355 ;
        RECT 633.255 123.975 636.555 124.355 ;
        RECT 637.255 123.975 638.615 124.355 ;
        RECT 640.590 123.975 642.055 124.355 ;
        RECT 642.755 123.975 646.055 124.355 ;
        RECT 646.755 123.975 650.055 124.355 ;
        RECT 650.755 123.975 651.935 124.355 ;
        RECT 665.650 123.950 666.955 124.330 ;
        RECT 671.655 123.950 674.955 124.330 ;
        RECT 675.655 123.950 677.015 124.330 ;
        RECT 678.990 123.950 680.455 124.330 ;
        RECT 681.155 123.950 684.455 124.330 ;
        RECT 689.155 123.950 690.335 124.330 ;
        RECT 628.715 123.630 629.095 123.665 ;
        RECT 610.750 123.145 611.130 123.525 ;
        RECT 613.155 123.160 614.935 123.450 ;
        RECT 616.410 123.250 617.600 123.535 ;
        RECT 620.530 123.130 621.840 123.450 ;
        RECT 628.450 123.320 631.460 123.630 ;
        RECT 628.715 123.285 629.095 123.320 ;
        RECT 632.715 123.285 633.805 123.665 ;
        RECT 636.715 123.660 637.095 123.665 ;
        RECT 634.235 123.295 637.100 123.660 ;
        RECT 642.215 123.640 642.595 123.665 ;
        RECT 642.200 123.320 644.345 123.640 ;
        RECT 636.715 123.285 637.095 123.295 ;
        RECT 642.215 123.285 642.595 123.320 ;
        RECT 645.260 123.285 646.595 123.665 ;
        RECT 650.215 123.645 650.595 123.665 ;
        RECT 647.750 123.325 650.660 123.645 ;
        RECT 667.115 123.605 667.495 123.640 ;
        RECT 650.215 123.285 650.595 123.325 ;
        RECT 666.850 123.295 669.860 123.605 ;
        RECT 667.115 123.260 667.495 123.295 ;
        RECT 671.115 123.260 672.205 123.640 ;
        RECT 675.115 123.635 675.495 123.640 ;
        RECT 672.635 123.270 675.500 123.635 ;
        RECT 680.615 123.615 680.995 123.640 ;
        RECT 680.600 123.295 682.745 123.615 ;
        RECT 675.115 123.260 675.495 123.270 ;
        RECT 680.615 123.260 680.995 123.295 ;
        RECT 683.660 123.260 684.995 123.640 ;
        RECT 688.615 123.620 688.995 123.640 ;
        RECT 686.150 123.300 689.060 123.620 ;
        RECT 688.615 123.260 688.995 123.300 ;
        RECT 693.245 123.120 693.625 123.500 ;
        RECT 695.650 123.135 697.430 123.425 ;
        RECT 698.905 123.225 700.095 123.510 ;
        RECT 703.025 123.105 704.335 123.425 ;
        RECT 611.885 122.545 612.265 122.925 ;
        RECT 615.630 122.585 616.010 122.965 ;
        RECT 618.340 122.575 618.720 122.955 ;
        RECT 619.750 122.420 622.930 122.740 ;
        RECT 694.380 122.520 694.760 122.900 ;
        RECT 698.125 122.560 698.505 122.940 ;
        RECT 700.835 122.550 701.215 122.930 ;
        RECT 702.245 122.395 705.425 122.715 ;
        RECT 627.065 121.975 628.555 122.355 ;
        RECT 629.255 121.975 630.540 122.355 ;
        RECT 648.570 121.975 650.055 122.355 ;
        RECT 650.755 121.975 651.830 122.355 ;
        RECT 665.465 121.950 666.955 122.330 ;
        RECT 689.155 121.950 690.230 122.330 ;
        RECT 628.715 121.285 629.805 121.665 ;
        RECT 630.760 121.295 632.280 121.655 ;
        RECT 633.200 121.290 646.050 121.625 ;
        RECT 650.215 121.620 650.595 121.665 ;
        RECT 649.480 121.320 650.790 121.620 ;
        RECT 650.215 121.285 650.595 121.320 ;
        RECT 667.115 121.260 668.205 121.640 ;
        RECT 669.160 121.270 670.680 121.630 ;
        RECT 671.600 121.265 684.450 121.600 ;
        RECT 688.615 121.595 688.995 121.640 ;
        RECT 687.880 121.295 689.190 121.595 ;
        RECT 688.615 121.260 688.995 121.295 ;
        RECT 625.570 120.765 658.650 120.775 ;
        RECT 625.570 120.425 690.625 120.765 ;
        RECT 657.675 120.400 690.625 120.425 ;
        RECT 692.420 120.390 696.680 120.745 ;
        RECT 609.680 119.830 613.775 119.835 ;
        RECT 593.100 119.825 598.315 119.830 ;
        RECT 608.560 119.825 613.775 119.830 ;
        RECT 624.020 119.825 664.270 119.830 ;
        RECT 593.100 119.805 664.270 119.825 ;
        RECT 690.625 119.805 696.270 119.810 ;
        RECT 706.885 119.805 707.265 125.635 ;
        RECT 715.765 125.585 720.265 125.895 ;
        RECT 792.185 125.660 796.315 125.960 ;
        RECT 711.725 125.035 718.115 125.325 ;
        RECT 711.140 124.455 727.160 124.790 ;
        RECT 775.945 124.555 781.860 124.890 ;
        RECT 779.215 124.535 781.860 124.555 ;
        RECT 710.490 123.870 713.410 124.170 ;
        RECT 716.955 123.855 720.325 124.155 ;
        RECT 756.540 123.915 759.840 124.295 ;
        RECT 760.540 123.915 763.840 124.295 ;
        RECT 770.040 123.915 773.340 124.295 ;
        RECT 774.040 123.915 777.340 124.295 ;
        RECT 708.705 123.120 709.085 123.500 ;
        RECT 711.110 123.135 712.890 123.425 ;
        RECT 714.365 123.225 715.555 123.510 ;
        RECT 718.485 123.105 719.795 123.425 ;
        RECT 709.840 122.520 710.220 122.900 ;
        RECT 713.585 122.560 713.965 122.940 ;
        RECT 716.295 122.550 716.675 122.930 ;
        RECT 717.705 122.395 720.885 122.715 ;
        RECT 756.540 121.915 757.825 122.295 ;
        RECT 775.855 121.915 777.340 122.295 ;
        RECT 707.985 121.310 712.135 121.580 ;
        RECT 758.045 121.235 759.565 121.595 ;
        RECT 789.810 119.830 790.190 125.660 ;
        RECT 798.690 125.610 803.190 125.920 ;
        RECT 807.645 125.660 811.775 125.960 ;
        RECT 794.650 125.060 801.040 125.350 ;
        RECT 794.065 124.480 804.720 124.815 ;
        RECT 793.415 123.895 796.335 124.195 ;
        RECT 799.880 123.880 803.250 124.180 ;
        RECT 791.630 123.145 792.010 123.525 ;
        RECT 794.035 123.160 795.815 123.450 ;
        RECT 797.290 123.250 798.480 123.535 ;
        RECT 801.410 123.130 802.720 123.450 ;
        RECT 792.765 122.545 793.145 122.925 ;
        RECT 796.510 122.585 796.890 122.965 ;
        RECT 799.220 122.575 799.600 122.955 ;
        RECT 800.630 122.420 803.810 122.740 ;
        RECT 790.560 119.830 794.655 119.835 ;
        RECT 805.270 119.830 805.650 125.660 ;
        RECT 814.150 125.610 818.650 125.920 ;
        RECT 905.600 125.635 909.730 125.935 ;
        RECT 821.380 125.425 857.290 125.450 ;
        RECT 810.110 125.060 816.500 125.350 ;
        RECT 821.380 125.180 888.385 125.425 ;
        RECT 856.640 125.155 888.385 125.180 ;
        RECT 892.605 125.035 898.995 125.325 ;
        RECT 809.525 124.480 820.030 124.815 ;
        RECT 845.000 124.615 855.550 124.950 ;
        RECT 892.020 124.455 902.500 124.790 ;
        RECT 808.875 123.895 811.795 124.195 ;
        RECT 815.340 123.880 818.710 124.180 ;
        RECT 823.590 123.975 824.895 124.355 ;
        RECT 825.595 123.975 828.895 124.355 ;
        RECT 829.595 123.975 832.895 124.355 ;
        RECT 833.595 123.975 834.955 124.355 ;
        RECT 836.930 123.975 838.395 124.355 ;
        RECT 839.095 123.975 842.395 124.355 ;
        RECT 843.095 123.975 846.395 124.355 ;
        RECT 847.095 123.975 848.275 124.355 ;
        RECT 861.990 123.950 863.295 124.330 ;
        RECT 867.995 123.950 871.295 124.330 ;
        RECT 871.995 123.950 873.355 124.330 ;
        RECT 875.330 123.950 876.795 124.330 ;
        RECT 877.495 123.950 880.795 124.330 ;
        RECT 885.495 123.950 886.675 124.330 ;
        RECT 825.055 123.630 825.435 123.665 ;
        RECT 807.090 123.145 807.470 123.525 ;
        RECT 809.495 123.160 811.275 123.450 ;
        RECT 812.750 123.250 813.940 123.535 ;
        RECT 816.870 123.130 818.180 123.450 ;
        RECT 824.790 123.320 827.800 123.630 ;
        RECT 825.055 123.285 825.435 123.320 ;
        RECT 829.055 123.285 830.145 123.665 ;
        RECT 833.055 123.660 833.435 123.665 ;
        RECT 830.575 123.295 833.440 123.660 ;
        RECT 838.555 123.640 838.935 123.665 ;
        RECT 838.540 123.320 840.685 123.640 ;
        RECT 833.055 123.285 833.435 123.295 ;
        RECT 838.555 123.285 838.935 123.320 ;
        RECT 841.600 123.285 842.935 123.665 ;
        RECT 846.555 123.645 846.935 123.665 ;
        RECT 844.090 123.325 847.000 123.645 ;
        RECT 863.455 123.605 863.835 123.640 ;
        RECT 846.555 123.285 846.935 123.325 ;
        RECT 863.190 123.295 866.200 123.605 ;
        RECT 863.455 123.260 863.835 123.295 ;
        RECT 867.455 123.260 868.545 123.640 ;
        RECT 871.455 123.635 871.835 123.640 ;
        RECT 868.975 123.270 871.840 123.635 ;
        RECT 876.955 123.615 877.335 123.640 ;
        RECT 876.940 123.295 879.085 123.615 ;
        RECT 871.455 123.260 871.835 123.270 ;
        RECT 876.955 123.260 877.335 123.295 ;
        RECT 880.000 123.260 881.335 123.640 ;
        RECT 884.955 123.620 885.335 123.640 ;
        RECT 882.490 123.300 885.400 123.620 ;
        RECT 884.955 123.260 885.335 123.300 ;
        RECT 889.585 123.120 889.965 123.500 ;
        RECT 891.990 123.135 893.770 123.425 ;
        RECT 895.245 123.225 896.435 123.510 ;
        RECT 899.365 123.105 900.675 123.425 ;
        RECT 808.225 122.545 808.605 122.925 ;
        RECT 811.970 122.585 812.350 122.965 ;
        RECT 814.680 122.575 815.060 122.955 ;
        RECT 816.090 122.420 819.270 122.740 ;
        RECT 890.720 122.520 891.100 122.900 ;
        RECT 894.465 122.560 894.845 122.940 ;
        RECT 897.175 122.550 897.555 122.930 ;
        RECT 898.585 122.395 901.765 122.715 ;
        RECT 823.405 121.975 824.895 122.355 ;
        RECT 825.595 121.975 826.880 122.355 ;
        RECT 844.910 121.975 846.395 122.355 ;
        RECT 847.095 121.975 848.170 122.355 ;
        RECT 861.805 121.950 863.295 122.330 ;
        RECT 885.495 121.950 886.570 122.330 ;
        RECT 825.055 121.285 826.145 121.665 ;
        RECT 827.100 121.295 828.620 121.655 ;
        RECT 829.540 121.290 842.390 121.625 ;
        RECT 846.555 121.620 846.935 121.665 ;
        RECT 845.820 121.320 847.130 121.620 ;
        RECT 846.555 121.285 846.935 121.320 ;
        RECT 863.455 121.260 864.545 121.640 ;
        RECT 865.500 121.270 867.020 121.630 ;
        RECT 867.940 121.265 880.790 121.600 ;
        RECT 884.955 121.595 885.335 121.640 ;
        RECT 884.220 121.295 885.530 121.595 ;
        RECT 884.955 121.260 885.335 121.295 ;
        RECT 821.910 120.765 854.990 120.775 ;
        RECT 821.910 120.425 886.965 120.765 ;
        RECT 854.015 120.400 886.965 120.425 ;
        RECT 888.760 120.390 893.020 120.745 ;
        RECT 806.020 119.830 810.115 119.835 ;
        RECT 789.440 119.825 794.655 119.830 ;
        RECT 804.900 119.825 810.115 119.830 ;
        RECT 820.360 119.825 860.610 119.830 ;
        RECT 707.635 119.805 711.730 119.810 ;
        RECT 593.100 119.800 696.270 119.805 ;
        RECT 706.515 119.800 711.730 119.805 ;
        RECT 789.440 119.805 860.610 119.825 ;
        RECT 886.965 119.805 892.610 119.810 ;
        RECT 903.225 119.805 903.605 125.635 ;
        RECT 912.105 125.585 916.605 125.895 ;
        RECT 988.525 125.660 992.655 125.960 ;
        RECT 908.065 125.035 914.455 125.325 ;
        RECT 907.480 124.455 923.500 124.790 ;
        RECT 972.330 124.540 978.245 124.875 ;
        RECT 975.600 124.520 978.245 124.540 ;
        RECT 906.830 123.870 909.750 124.170 ;
        RECT 913.295 123.855 916.665 124.155 ;
        RECT 952.925 123.900 956.225 124.280 ;
        RECT 956.925 123.900 960.225 124.280 ;
        RECT 966.425 123.900 969.725 124.280 ;
        RECT 970.425 123.900 973.725 124.280 ;
        RECT 905.045 123.120 905.425 123.500 ;
        RECT 907.450 123.135 909.230 123.425 ;
        RECT 910.705 123.225 911.895 123.510 ;
        RECT 914.825 123.105 916.135 123.425 ;
        RECT 906.180 122.520 906.560 122.900 ;
        RECT 909.925 122.560 910.305 122.940 ;
        RECT 912.635 122.550 913.015 122.930 ;
        RECT 914.045 122.395 917.225 122.715 ;
        RECT 952.925 121.900 954.210 122.280 ;
        RECT 972.240 121.900 973.725 122.280 ;
        RECT 904.325 121.310 908.475 121.580 ;
        RECT 954.430 121.220 955.950 121.580 ;
        RECT 986.150 119.830 986.530 125.660 ;
        RECT 995.030 125.610 999.530 125.920 ;
        RECT 1003.985 125.660 1008.115 125.960 ;
        RECT 990.990 125.060 997.380 125.350 ;
        RECT 990.405 124.480 1001.060 124.815 ;
        RECT 989.755 123.895 992.675 124.195 ;
        RECT 996.220 123.880 999.590 124.180 ;
        RECT 987.970 123.145 988.350 123.525 ;
        RECT 990.375 123.160 992.155 123.450 ;
        RECT 993.630 123.250 994.820 123.535 ;
        RECT 997.750 123.130 999.060 123.450 ;
        RECT 989.105 122.545 989.485 122.925 ;
        RECT 992.850 122.585 993.230 122.965 ;
        RECT 995.560 122.575 995.940 122.955 ;
        RECT 996.970 122.420 1000.150 122.740 ;
        RECT 986.900 119.830 990.995 119.835 ;
        RECT 1001.610 119.830 1001.990 125.660 ;
        RECT 1010.490 125.610 1014.990 125.920 ;
        RECT 1101.940 125.635 1106.070 125.935 ;
        RECT 1017.720 125.425 1053.630 125.450 ;
        RECT 1006.450 125.060 1012.840 125.350 ;
        RECT 1017.720 125.180 1084.725 125.425 ;
        RECT 1052.980 125.155 1084.725 125.180 ;
        RECT 1088.945 125.035 1095.335 125.325 ;
        RECT 1005.865 124.480 1016.370 124.815 ;
        RECT 1041.340 124.615 1051.890 124.950 ;
        RECT 1088.360 124.455 1098.840 124.790 ;
        RECT 1005.215 123.895 1008.135 124.195 ;
        RECT 1011.680 123.880 1015.050 124.180 ;
        RECT 1019.930 123.975 1021.235 124.355 ;
        RECT 1021.935 123.975 1025.235 124.355 ;
        RECT 1025.935 123.975 1029.235 124.355 ;
        RECT 1029.935 123.975 1031.295 124.355 ;
        RECT 1033.270 123.975 1034.735 124.355 ;
        RECT 1035.435 123.975 1038.735 124.355 ;
        RECT 1039.435 123.975 1042.735 124.355 ;
        RECT 1043.435 123.975 1044.615 124.355 ;
        RECT 1058.330 123.950 1059.635 124.330 ;
        RECT 1064.335 123.950 1067.635 124.330 ;
        RECT 1068.335 123.950 1069.695 124.330 ;
        RECT 1071.670 123.950 1073.135 124.330 ;
        RECT 1073.835 123.950 1077.135 124.330 ;
        RECT 1081.835 123.950 1083.015 124.330 ;
        RECT 1021.395 123.630 1021.775 123.665 ;
        RECT 1003.430 123.145 1003.810 123.525 ;
        RECT 1005.835 123.160 1007.615 123.450 ;
        RECT 1009.090 123.250 1010.280 123.535 ;
        RECT 1013.210 123.130 1014.520 123.450 ;
        RECT 1021.130 123.320 1024.140 123.630 ;
        RECT 1021.395 123.285 1021.775 123.320 ;
        RECT 1025.395 123.285 1026.485 123.665 ;
        RECT 1029.395 123.660 1029.775 123.665 ;
        RECT 1026.915 123.295 1029.780 123.660 ;
        RECT 1034.895 123.640 1035.275 123.665 ;
        RECT 1034.880 123.320 1037.025 123.640 ;
        RECT 1029.395 123.285 1029.775 123.295 ;
        RECT 1034.895 123.285 1035.275 123.320 ;
        RECT 1037.940 123.285 1039.275 123.665 ;
        RECT 1042.895 123.645 1043.275 123.665 ;
        RECT 1040.430 123.325 1043.340 123.645 ;
        RECT 1059.795 123.605 1060.175 123.640 ;
        RECT 1042.895 123.285 1043.275 123.325 ;
        RECT 1059.530 123.295 1062.540 123.605 ;
        RECT 1059.795 123.260 1060.175 123.295 ;
        RECT 1063.795 123.260 1064.885 123.640 ;
        RECT 1067.795 123.635 1068.175 123.640 ;
        RECT 1065.315 123.270 1068.180 123.635 ;
        RECT 1073.295 123.615 1073.675 123.640 ;
        RECT 1073.280 123.295 1075.425 123.615 ;
        RECT 1067.795 123.260 1068.175 123.270 ;
        RECT 1073.295 123.260 1073.675 123.295 ;
        RECT 1076.340 123.260 1077.675 123.640 ;
        RECT 1081.295 123.620 1081.675 123.640 ;
        RECT 1078.830 123.300 1081.740 123.620 ;
        RECT 1081.295 123.260 1081.675 123.300 ;
        RECT 1085.925 123.120 1086.305 123.500 ;
        RECT 1088.330 123.135 1090.110 123.425 ;
        RECT 1091.585 123.225 1092.775 123.510 ;
        RECT 1095.705 123.105 1097.015 123.425 ;
        RECT 1004.565 122.545 1004.945 122.925 ;
        RECT 1008.310 122.585 1008.690 122.965 ;
        RECT 1011.020 122.575 1011.400 122.955 ;
        RECT 1012.430 122.420 1015.610 122.740 ;
        RECT 1087.060 122.520 1087.440 122.900 ;
        RECT 1090.805 122.560 1091.185 122.940 ;
        RECT 1093.515 122.550 1093.895 122.930 ;
        RECT 1094.925 122.395 1098.105 122.715 ;
        RECT 1019.745 121.975 1021.235 122.355 ;
        RECT 1021.935 121.975 1023.220 122.355 ;
        RECT 1041.250 121.975 1042.735 122.355 ;
        RECT 1043.435 121.975 1044.510 122.355 ;
        RECT 1058.145 121.950 1059.635 122.330 ;
        RECT 1081.835 121.950 1082.910 122.330 ;
        RECT 1021.395 121.285 1022.485 121.665 ;
        RECT 1023.440 121.295 1024.960 121.655 ;
        RECT 1025.880 121.290 1038.730 121.625 ;
        RECT 1042.895 121.620 1043.275 121.665 ;
        RECT 1042.160 121.320 1043.470 121.620 ;
        RECT 1042.895 121.285 1043.275 121.320 ;
        RECT 1059.795 121.260 1060.885 121.640 ;
        RECT 1061.840 121.270 1063.360 121.630 ;
        RECT 1064.280 121.265 1077.130 121.600 ;
        RECT 1081.295 121.595 1081.675 121.640 ;
        RECT 1080.560 121.295 1081.870 121.595 ;
        RECT 1081.295 121.260 1081.675 121.295 ;
        RECT 1018.250 120.765 1051.330 120.775 ;
        RECT 1018.250 120.425 1083.305 120.765 ;
        RECT 1050.355 120.400 1083.305 120.425 ;
        RECT 1085.100 120.390 1089.360 120.745 ;
        RECT 1002.360 119.830 1006.455 119.835 ;
        RECT 985.780 119.825 990.995 119.830 ;
        RECT 1001.240 119.825 1006.455 119.830 ;
        RECT 1016.700 119.825 1056.950 119.830 ;
        RECT 903.975 119.805 908.070 119.810 ;
        RECT 789.440 119.800 892.610 119.805 ;
        RECT 902.855 119.800 908.070 119.805 ;
        RECT 985.780 119.805 1056.950 119.825 ;
        RECT 1083.305 119.805 1088.950 119.810 ;
        RECT 1099.565 119.805 1099.945 125.635 ;
        RECT 1108.445 125.585 1112.945 125.895 ;
        RECT 1184.865 125.660 1188.995 125.960 ;
        RECT 1104.405 125.035 1110.795 125.325 ;
        RECT 1103.820 124.455 1119.840 124.790 ;
        RECT 1168.655 124.545 1174.570 124.880 ;
        RECT 1171.925 124.525 1174.570 124.545 ;
        RECT 1103.170 123.870 1106.090 124.170 ;
        RECT 1109.635 123.855 1113.005 124.155 ;
        RECT 1149.250 123.905 1152.550 124.285 ;
        RECT 1153.250 123.905 1156.550 124.285 ;
        RECT 1162.750 123.905 1166.050 124.285 ;
        RECT 1166.750 123.905 1170.050 124.285 ;
        RECT 1101.385 123.120 1101.765 123.500 ;
        RECT 1103.790 123.135 1105.570 123.425 ;
        RECT 1107.045 123.225 1108.235 123.510 ;
        RECT 1111.165 123.105 1112.475 123.425 ;
        RECT 1102.520 122.520 1102.900 122.900 ;
        RECT 1106.265 122.560 1106.645 122.940 ;
        RECT 1108.975 122.550 1109.355 122.930 ;
        RECT 1110.385 122.395 1113.565 122.715 ;
        RECT 1149.250 121.905 1150.535 122.285 ;
        RECT 1168.565 121.905 1170.050 122.285 ;
        RECT 1100.665 121.310 1104.815 121.580 ;
        RECT 1150.755 121.225 1152.275 121.585 ;
        RECT 1182.490 119.830 1182.870 125.660 ;
        RECT 1191.370 125.610 1195.870 125.920 ;
        RECT 1200.325 125.660 1204.455 125.960 ;
        RECT 1187.330 125.060 1193.720 125.350 ;
        RECT 1186.745 124.480 1197.400 124.815 ;
        RECT 1186.095 123.895 1189.015 124.195 ;
        RECT 1192.560 123.880 1195.930 124.180 ;
        RECT 1184.310 123.145 1184.690 123.525 ;
        RECT 1186.715 123.160 1188.495 123.450 ;
        RECT 1189.970 123.250 1191.160 123.535 ;
        RECT 1194.090 123.130 1195.400 123.450 ;
        RECT 1185.445 122.545 1185.825 122.925 ;
        RECT 1189.190 122.585 1189.570 122.965 ;
        RECT 1191.900 122.575 1192.280 122.955 ;
        RECT 1193.310 122.420 1196.490 122.740 ;
        RECT 1183.240 119.830 1187.335 119.835 ;
        RECT 1197.950 119.830 1198.330 125.660 ;
        RECT 1206.830 125.610 1211.330 125.920 ;
        RECT 1282.820 125.635 1286.950 125.935 ;
        RECT 1289.325 125.585 1293.825 125.895 ;
        RECT 1298.280 125.635 1302.410 125.935 ;
        RECT 1214.060 125.425 1249.970 125.450 ;
        RECT 1202.790 125.060 1209.180 125.350 ;
        RECT 1214.060 125.180 1281.065 125.425 ;
        RECT 1249.320 125.155 1281.065 125.180 ;
        RECT 1285.285 125.035 1291.675 125.325 ;
        RECT 1202.205 124.480 1212.710 124.815 ;
        RECT 1237.680 124.615 1248.230 124.950 ;
        RECT 1276.080 124.590 1280.025 124.925 ;
        RECT 1284.700 124.455 1295.180 124.790 ;
        RECT 1201.555 123.895 1204.475 124.195 ;
        RECT 1208.020 123.880 1211.390 124.180 ;
        RECT 1216.270 123.975 1217.575 124.355 ;
        RECT 1218.275 123.975 1221.575 124.355 ;
        RECT 1222.275 123.975 1225.575 124.355 ;
        RECT 1226.275 123.975 1227.635 124.355 ;
        RECT 1229.610 123.975 1231.075 124.355 ;
        RECT 1231.775 123.975 1235.075 124.355 ;
        RECT 1235.775 123.975 1239.075 124.355 ;
        RECT 1239.775 123.975 1240.955 124.355 ;
        RECT 1254.670 123.950 1255.975 124.330 ;
        RECT 1256.675 123.950 1259.975 124.330 ;
        RECT 1260.675 123.950 1263.975 124.330 ;
        RECT 1264.675 123.950 1266.035 124.330 ;
        RECT 1268.010 123.950 1269.475 124.330 ;
        RECT 1270.175 123.950 1273.475 124.330 ;
        RECT 1274.175 123.950 1277.475 124.330 ;
        RECT 1278.175 123.950 1279.355 124.330 ;
        RECT 1284.050 123.870 1286.970 124.170 ;
        RECT 1290.515 123.855 1293.885 124.155 ;
        RECT 1217.735 123.630 1218.115 123.665 ;
        RECT 1199.770 123.145 1200.150 123.525 ;
        RECT 1202.175 123.160 1203.955 123.450 ;
        RECT 1205.430 123.250 1206.620 123.535 ;
        RECT 1209.550 123.130 1210.860 123.450 ;
        RECT 1217.470 123.320 1220.480 123.630 ;
        RECT 1217.735 123.285 1218.115 123.320 ;
        RECT 1221.735 123.285 1222.825 123.665 ;
        RECT 1225.735 123.660 1226.115 123.665 ;
        RECT 1223.255 123.295 1226.120 123.660 ;
        RECT 1231.235 123.640 1231.615 123.665 ;
        RECT 1231.220 123.320 1233.365 123.640 ;
        RECT 1225.735 123.285 1226.115 123.295 ;
        RECT 1231.235 123.285 1231.615 123.320 ;
        RECT 1234.280 123.285 1235.615 123.665 ;
        RECT 1239.235 123.645 1239.615 123.665 ;
        RECT 1236.770 123.325 1239.680 123.645 ;
        RECT 1256.135 123.605 1256.515 123.640 ;
        RECT 1239.235 123.285 1239.615 123.325 ;
        RECT 1255.870 123.295 1258.880 123.605 ;
        RECT 1256.135 123.260 1256.515 123.295 ;
        RECT 1260.135 123.260 1261.225 123.640 ;
        RECT 1264.135 123.635 1264.515 123.640 ;
        RECT 1261.655 123.270 1264.520 123.635 ;
        RECT 1269.635 123.615 1270.015 123.640 ;
        RECT 1269.620 123.295 1271.765 123.615 ;
        RECT 1264.135 123.260 1264.515 123.270 ;
        RECT 1269.635 123.260 1270.015 123.295 ;
        RECT 1272.680 123.260 1274.015 123.640 ;
        RECT 1277.635 123.620 1278.015 123.640 ;
        RECT 1275.170 123.300 1278.080 123.620 ;
        RECT 1277.635 123.260 1278.015 123.300 ;
        RECT 1282.265 123.120 1282.645 123.500 ;
        RECT 1284.670 123.135 1286.450 123.425 ;
        RECT 1287.925 123.225 1289.115 123.510 ;
        RECT 1292.045 123.105 1293.355 123.425 ;
        RECT 1200.905 122.545 1201.285 122.925 ;
        RECT 1204.650 122.585 1205.030 122.965 ;
        RECT 1207.360 122.575 1207.740 122.955 ;
        RECT 1208.770 122.420 1211.950 122.740 ;
        RECT 1283.400 122.520 1283.780 122.900 ;
        RECT 1287.145 122.560 1287.525 122.940 ;
        RECT 1289.855 122.550 1290.235 122.930 ;
        RECT 1291.265 122.395 1294.445 122.715 ;
        RECT 1216.085 121.975 1217.575 122.355 ;
        RECT 1218.275 121.975 1219.560 122.355 ;
        RECT 1237.590 121.975 1239.075 122.355 ;
        RECT 1239.775 121.975 1240.850 122.355 ;
        RECT 1254.485 121.950 1255.975 122.330 ;
        RECT 1256.675 121.950 1257.960 122.330 ;
        RECT 1275.990 121.950 1277.475 122.330 ;
        RECT 1278.175 121.950 1279.250 122.330 ;
        RECT 1217.735 121.285 1218.825 121.665 ;
        RECT 1219.780 121.295 1221.300 121.655 ;
        RECT 1222.220 121.290 1235.070 121.625 ;
        RECT 1239.235 121.620 1239.615 121.665 ;
        RECT 1238.500 121.320 1239.810 121.620 ;
        RECT 1239.235 121.285 1239.615 121.320 ;
        RECT 1256.135 121.260 1257.225 121.640 ;
        RECT 1258.180 121.270 1259.700 121.630 ;
        RECT 1260.620 121.265 1273.470 121.600 ;
        RECT 1277.635 121.595 1278.015 121.640 ;
        RECT 1276.900 121.295 1278.210 121.595 ;
        RECT 1277.635 121.260 1278.015 121.295 ;
        RECT 1214.590 120.765 1247.670 120.775 ;
        RECT 1214.590 120.425 1279.645 120.765 ;
        RECT 1246.695 120.400 1279.645 120.425 ;
        RECT 1281.440 120.390 1285.700 120.745 ;
        RECT 1198.700 119.830 1202.795 119.835 ;
        RECT 1182.120 119.825 1187.335 119.830 ;
        RECT 1197.580 119.825 1202.795 119.830 ;
        RECT 1213.040 119.825 1253.290 119.830 ;
        RECT 1100.315 119.805 1104.410 119.810 ;
        RECT 985.780 119.800 1088.950 119.805 ;
        RECT 1099.195 119.800 1104.410 119.805 ;
        RECT 1182.120 119.805 1253.290 119.825 ;
        RECT 1279.645 119.805 1285.290 119.810 ;
        RECT 1295.905 119.805 1296.285 125.635 ;
        RECT 1304.785 125.585 1309.285 125.895 ;
        RECT 1300.745 125.035 1307.135 125.325 ;
        RECT 1299.510 123.870 1302.430 124.170 ;
        RECT 1305.975 123.855 1309.345 124.155 ;
        RECT 1297.725 123.120 1298.105 123.500 ;
        RECT 1303.385 123.225 1304.575 123.510 ;
        RECT 1302.605 122.560 1302.985 122.940 ;
        RECT 1306.725 122.395 1309.905 122.715 ;
        RECT 1297.005 121.310 1301.155 121.580 ;
        RECT 1296.655 119.805 1300.750 119.810 ;
        RECT 1182.120 119.800 1285.290 119.805 ;
        RECT 1295.535 119.800 1300.750 119.805 ;
        RECT 511.260 119.770 515.355 119.775 ;
        RECT 396.725 119.765 499.895 119.770 ;
        RECT 510.140 119.765 515.355 119.770 ;
        RECT 271.195 118.920 328.770 118.945 ;
        RECT 360.170 118.820 386.825 119.720 ;
        RECT 396.725 118.895 525.170 119.765 ;
        RECT 467.595 118.870 525.170 118.895 ;
        RECT 556.490 118.865 583.145 119.765 ;
        RECT 593.100 118.930 721.545 119.800 ;
        RECT 663.970 118.905 721.545 118.930 ;
        RECT 752.855 118.870 779.510 119.770 ;
        RECT 789.440 118.930 917.885 119.800 ;
        RECT 860.310 118.905 917.885 118.930 ;
        RECT 949.240 118.855 975.895 119.755 ;
        RECT 985.780 118.930 1114.225 119.800 ;
        RECT 1056.650 118.905 1114.225 118.930 ;
        RECT 1145.565 118.860 1172.220 119.760 ;
        RECT 1182.120 118.930 1310.565 119.800 ;
        RECT 1252.990 118.905 1310.565 118.930 ;
        RECT 76.050 115.030 132.405 115.050 ;
        RECT 272.415 115.030 328.770 115.050 ;
        RECT -81.565 114.025 -56.130 114.925 ;
        RECT -31.240 114.105 -5.805 115.005 ;
        RECT 3.765 114.150 132.405 115.030 ;
        RECT 3.765 114.130 76.155 114.150 ;
        RECT -79.080 111.845 -77.880 112.225 ;
        RECT -76.125 111.630 -73.850 112.140 ;
        RECT -71.225 111.630 -68.925 112.140 ;
        RECT -66.630 111.630 -64.350 112.140 ;
        RECT -59.555 111.945 -58.320 112.325 ;
        RECT -28.755 111.925 -27.555 112.305 ;
        RECT -25.800 111.710 -23.525 112.220 ;
        RECT -20.900 111.710 -18.600 112.220 ;
        RECT -16.305 111.710 -14.025 112.220 ;
        RECT -9.230 112.025 -7.995 112.405 ;
        RECT -79.080 109.545 -75.820 109.925 ;
        RECT -75.080 109.545 -71.820 109.925 ;
        RECT -65.580 109.545 -62.320 109.925 ;
        RECT -61.580 109.545 -58.320 109.925 ;
        RECT -28.755 109.625 -25.495 110.005 ;
        RECT -24.755 109.625 -21.495 110.005 ;
        RECT -15.255 109.625 -11.995 110.005 ;
        RECT -11.255 109.625 -7.995 110.005 ;
        RECT -78.415 107.960 -56.130 107.970 ;
        RECT -78.415 107.630 -54.590 107.960 ;
        RECT -28.090 107.710 -1.795 108.050 ;
        RECT -56.350 107.610 -54.590 107.630 ;
        RECT 4.135 106.970 4.515 114.130 ;
        RECT 5.965 109.915 9.340 110.315 ;
        RECT 9.710 109.675 10.090 110.055 ;
        RECT 12.425 109.715 12.805 110.095 ;
        RECT 16.610 109.665 16.990 110.045 ;
        RECT 7.035 109.250 8.775 109.540 ;
        RECT 10.825 109.200 12.025 109.490 ;
        RECT 13.535 109.170 16.145 109.595 ;
        RECT 17.745 109.265 18.125 109.645 ;
        RECT 5.280 108.490 18.845 108.805 ;
        RECT 5.275 107.745 18.835 108.045 ;
        RECT 5.295 107.030 12.020 107.330 ;
        RECT 15.720 106.730 18.825 107.005 ;
        RECT 19.595 106.970 19.975 114.130 ;
        RECT 73.035 113.145 101.810 113.165 ;
        RECT 36.235 112.880 101.810 113.145 ;
        RECT 36.235 112.860 73.785 112.880 ;
        RECT 103.480 112.860 110.185 113.160 ;
        RECT 37.745 111.950 39.200 112.330 ;
        RECT 39.940 111.950 41.140 112.330 ;
        RECT 42.895 111.735 45.170 112.245 ;
        RECT 47.795 111.735 50.095 112.245 ;
        RECT 52.390 111.735 54.670 112.245 ;
        RECT 59.465 112.050 60.700 112.430 ;
        RECT 61.440 112.050 62.720 112.430 ;
        RECT 76.340 111.970 77.795 112.350 ;
        RECT 81.490 111.755 83.765 112.265 ;
        RECT 86.390 111.755 88.690 112.265 ;
        RECT 90.985 111.755 93.265 112.265 ;
        RECT 100.035 112.070 101.315 112.450 ;
        RECT 60.880 111.695 61.260 111.730 ;
        RECT 99.475 111.715 99.855 111.750 ;
        RECT 39.380 111.590 39.760 111.630 ;
        RECT 39.310 111.285 42.145 111.590 ;
        RECT 58.125 111.385 61.260 111.695 ;
        RECT 77.975 111.610 78.355 111.650 ;
        RECT 60.880 111.350 61.260 111.385 ;
        RECT 77.905 111.305 80.740 111.610 ;
        RECT 96.720 111.405 99.855 111.715 ;
        RECT 99.475 111.370 99.855 111.405 ;
        RECT 39.380 111.250 39.760 111.285 ;
        RECT 77.975 111.270 78.355 111.305 ;
        RECT 21.425 109.875 24.830 110.315 ;
        RECT 25.170 109.675 25.550 110.055 ;
        RECT 27.885 109.715 28.265 110.095 ;
        RECT 32.070 109.665 32.450 110.045 ;
        RECT 37.905 109.650 39.200 110.030 ;
        RECT 39.940 109.650 43.200 110.030 ;
        RECT 43.940 109.650 47.200 110.030 ;
        RECT 47.940 109.650 49.125 110.030 ;
        RECT 51.390 109.650 52.700 110.030 ;
        RECT 53.440 109.650 56.700 110.030 ;
        RECT 57.440 109.650 60.700 110.030 ;
        RECT 61.440 109.650 62.455 110.030 ;
        RECT 76.500 109.670 77.795 110.050 ;
        RECT 82.535 109.670 85.795 110.050 ;
        RECT 86.535 109.670 87.720 110.050 ;
        RECT 89.985 109.670 91.295 110.050 ;
        RECT 92.035 109.670 95.295 110.050 ;
        RECT 100.035 109.670 101.050 110.050 ;
        RECT 104.115 109.915 107.530 110.335 ;
        RECT 107.860 109.695 108.240 110.075 ;
        RECT 110.575 109.735 110.955 110.115 ;
        RECT 114.760 109.685 115.140 110.065 ;
        RECT 22.495 109.250 24.235 109.540 ;
        RECT 26.285 109.200 27.485 109.490 ;
        RECT 28.995 109.170 31.590 109.545 ;
        RECT 33.205 109.265 33.585 109.645 ;
        RECT 39.380 108.950 39.760 109.330 ;
        RECT 43.380 108.950 43.760 109.330 ;
        RECT 47.380 109.285 47.760 109.330 ;
        RECT 52.880 109.285 53.260 109.330 ;
        RECT 47.330 108.970 53.265 109.285 ;
        RECT 47.380 108.950 47.760 108.970 ;
        RECT 52.880 108.950 53.260 108.970 ;
        RECT 56.880 108.950 57.260 109.330 ;
        RECT 60.880 108.950 61.260 109.330 ;
        RECT 77.975 108.970 78.355 109.350 ;
        RECT 81.975 108.970 82.355 109.350 ;
        RECT 85.975 109.305 86.355 109.350 ;
        RECT 91.475 109.305 91.855 109.350 ;
        RECT 85.925 108.990 91.860 109.305 ;
        RECT 85.975 108.970 86.355 108.990 ;
        RECT 91.475 108.970 91.855 108.990 ;
        RECT 95.475 108.970 95.855 109.350 ;
        RECT 99.475 108.970 99.855 109.350 ;
        RECT 105.185 109.270 106.925 109.560 ;
        RECT 108.975 109.220 110.175 109.510 ;
        RECT 111.685 109.180 114.315 109.635 ;
        RECT 115.895 109.285 116.275 109.665 ;
        RECT 20.735 108.490 34.560 108.790 ;
        RECT 36.235 108.325 52.245 108.700 ;
        RECT 70.065 108.345 90.840 108.720 ;
        RECT 20.740 107.745 39.160 108.045 ;
        RECT 40.605 107.735 67.915 108.075 ;
        RECT 20.220 107.030 27.480 107.330 ;
        RECT 5.275 106.410 9.400 106.680 ;
        RECT 20.775 106.495 24.860 106.765 ;
        RECT 31.180 106.730 34.930 107.005 ;
        RECT 36.235 106.970 62.465 107.360 ;
        RECT 69.095 106.990 101.060 107.380 ;
        RECT 113.870 106.750 117.000 107.025 ;
        RECT 117.745 106.990 118.125 114.150 ;
        RECT 164.930 114.115 190.365 115.015 ;
        RECT 200.130 114.150 328.770 115.030 ;
        RECT 468.815 114.980 525.170 115.000 ;
        RECT 200.130 114.130 272.520 114.150 ;
        RECT 118.985 111.690 125.725 111.990 ;
        RECT 167.415 111.935 168.615 112.315 ;
        RECT 170.370 111.720 172.645 112.230 ;
        RECT 175.270 111.720 177.570 112.230 ;
        RECT 179.865 111.720 182.145 112.230 ;
        RECT 186.940 112.035 188.175 112.415 ;
        RECT 119.575 109.895 123.030 110.335 ;
        RECT 123.320 109.695 123.700 110.075 ;
        RECT 126.035 109.735 126.415 110.115 ;
        RECT 130.220 109.685 130.600 110.065 ;
        RECT 120.645 109.270 122.385 109.560 ;
        RECT 124.435 109.220 125.635 109.510 ;
        RECT 127.145 109.190 129.770 109.600 ;
        RECT 131.355 109.285 131.735 109.665 ;
        RECT 167.415 109.635 170.675 110.015 ;
        RECT 171.415 109.635 174.675 110.015 ;
        RECT 180.915 109.635 184.175 110.015 ;
        RECT 184.915 109.635 188.175 110.015 ;
        RECT 118.390 108.510 134.310 108.810 ;
        RECT 118.925 107.765 135.870 108.065 ;
        RECT 168.080 107.720 194.375 108.060 ;
        RECT 129.330 106.750 137.030 107.025 ;
        RECT 200.500 106.970 200.880 114.130 ;
        RECT 202.330 109.915 205.705 110.315 ;
        RECT 206.075 109.675 206.455 110.055 ;
        RECT 208.790 109.715 209.170 110.095 ;
        RECT 212.975 109.665 213.355 110.045 ;
        RECT 203.400 109.250 205.140 109.540 ;
        RECT 207.190 109.200 208.390 109.490 ;
        RECT 209.900 109.170 212.510 109.595 ;
        RECT 214.110 109.265 214.490 109.645 ;
        RECT 201.645 108.490 215.210 108.805 ;
        RECT 201.640 107.745 215.200 108.045 ;
        RECT 201.660 107.030 208.385 107.330 ;
        RECT 212.085 106.730 215.190 107.005 ;
        RECT 215.960 106.970 216.340 114.130 ;
        RECT 269.400 113.145 298.175 113.165 ;
        RECT 232.600 112.880 298.175 113.145 ;
        RECT 232.600 112.860 270.150 112.880 ;
        RECT 299.845 112.860 306.550 113.160 ;
        RECT 234.110 111.950 235.565 112.330 ;
        RECT 236.305 111.950 237.505 112.330 ;
        RECT 239.260 111.735 241.535 112.245 ;
        RECT 244.160 111.735 246.460 112.245 ;
        RECT 248.755 111.735 251.035 112.245 ;
        RECT 255.830 112.050 257.065 112.430 ;
        RECT 257.805 112.050 259.085 112.430 ;
        RECT 272.705 111.970 274.160 112.350 ;
        RECT 277.855 111.755 280.130 112.265 ;
        RECT 282.755 111.755 285.055 112.265 ;
        RECT 287.350 111.755 289.630 112.265 ;
        RECT 296.400 112.070 297.680 112.450 ;
        RECT 257.245 111.695 257.625 111.730 ;
        RECT 295.840 111.715 296.220 111.750 ;
        RECT 235.745 111.590 236.125 111.630 ;
        RECT 235.675 111.285 238.510 111.590 ;
        RECT 254.490 111.385 257.625 111.695 ;
        RECT 274.340 111.610 274.720 111.650 ;
        RECT 257.245 111.350 257.625 111.385 ;
        RECT 274.270 111.305 277.105 111.610 ;
        RECT 293.085 111.405 296.220 111.715 ;
        RECT 295.840 111.370 296.220 111.405 ;
        RECT 235.745 111.250 236.125 111.285 ;
        RECT 274.340 111.270 274.720 111.305 ;
        RECT 217.790 109.875 221.195 110.315 ;
        RECT 221.535 109.675 221.915 110.055 ;
        RECT 224.250 109.715 224.630 110.095 ;
        RECT 228.435 109.665 228.815 110.045 ;
        RECT 234.270 109.650 235.565 110.030 ;
        RECT 236.305 109.650 239.565 110.030 ;
        RECT 240.305 109.650 243.565 110.030 ;
        RECT 244.305 109.650 245.490 110.030 ;
        RECT 247.755 109.650 249.065 110.030 ;
        RECT 249.805 109.650 253.065 110.030 ;
        RECT 253.805 109.650 257.065 110.030 ;
        RECT 257.805 109.650 258.820 110.030 ;
        RECT 272.865 109.670 274.160 110.050 ;
        RECT 278.900 109.670 282.160 110.050 ;
        RECT 282.900 109.670 284.085 110.050 ;
        RECT 286.350 109.670 287.660 110.050 ;
        RECT 288.400 109.670 291.660 110.050 ;
        RECT 296.400 109.670 297.415 110.050 ;
        RECT 300.480 109.915 303.895 110.335 ;
        RECT 304.225 109.695 304.605 110.075 ;
        RECT 306.940 109.735 307.320 110.115 ;
        RECT 311.125 109.685 311.505 110.065 ;
        RECT 218.860 109.250 220.600 109.540 ;
        RECT 222.650 109.200 223.850 109.490 ;
        RECT 225.360 109.170 227.955 109.545 ;
        RECT 229.570 109.265 229.950 109.645 ;
        RECT 235.745 108.950 236.125 109.330 ;
        RECT 239.745 108.950 240.125 109.330 ;
        RECT 243.745 109.285 244.125 109.330 ;
        RECT 249.245 109.285 249.625 109.330 ;
        RECT 243.695 108.970 249.630 109.285 ;
        RECT 243.745 108.950 244.125 108.970 ;
        RECT 249.245 108.950 249.625 108.970 ;
        RECT 253.245 108.950 253.625 109.330 ;
        RECT 257.245 108.950 257.625 109.330 ;
        RECT 274.340 108.970 274.720 109.350 ;
        RECT 278.340 108.970 278.720 109.350 ;
        RECT 282.340 109.305 282.720 109.350 ;
        RECT 287.840 109.305 288.220 109.350 ;
        RECT 282.290 108.990 288.225 109.305 ;
        RECT 282.340 108.970 282.720 108.990 ;
        RECT 287.840 108.970 288.220 108.990 ;
        RECT 291.840 108.970 292.220 109.350 ;
        RECT 295.840 108.970 296.220 109.350 ;
        RECT 301.550 109.270 303.290 109.560 ;
        RECT 305.340 109.220 306.540 109.510 ;
        RECT 308.050 109.180 310.680 109.635 ;
        RECT 312.260 109.285 312.640 109.665 ;
        RECT 217.100 108.490 230.925 108.790 ;
        RECT 232.600 108.325 248.610 108.700 ;
        RECT 266.430 108.345 287.205 108.720 ;
        RECT 217.105 107.745 235.525 108.045 ;
        RECT 236.970 107.735 264.280 108.075 ;
        RECT 216.585 107.030 223.845 107.330 ;
        RECT 65.940 106.625 93.500 106.635 ;
        RECT 36.235 106.605 54.905 106.615 ;
        RECT 65.940 106.605 102.505 106.625 ;
        RECT 36.235 106.315 102.505 106.605 ;
        RECT 201.640 106.410 205.765 106.680 ;
        RECT 217.140 106.495 221.225 106.765 ;
        RECT 227.545 106.730 231.295 107.005 ;
        RECT 232.600 106.970 258.830 107.360 ;
        RECT 265.460 106.990 297.425 107.380 ;
        RECT 310.235 106.750 313.365 107.025 ;
        RECT 314.110 106.990 314.490 114.150 ;
        RECT 361.320 114.075 386.755 114.975 ;
        RECT 396.530 114.100 525.170 114.980 ;
        RECT 557.640 114.120 583.075 115.020 ;
        RECT 665.190 115.015 721.545 115.035 ;
        RECT 592.905 114.135 721.545 115.015 ;
        RECT 592.905 114.115 665.295 114.135 ;
        RECT 396.530 114.080 468.920 114.100 ;
        RECT 315.350 111.690 322.090 111.990 ;
        RECT 363.805 111.895 365.005 112.275 ;
        RECT 366.760 111.680 369.035 112.190 ;
        RECT 371.660 111.680 373.960 112.190 ;
        RECT 376.255 111.680 378.535 112.190 ;
        RECT 383.330 111.995 384.565 112.375 ;
        RECT 315.940 109.895 319.395 110.335 ;
        RECT 319.685 109.695 320.065 110.075 ;
        RECT 322.400 109.735 322.780 110.115 ;
        RECT 326.585 109.685 326.965 110.065 ;
        RECT 317.010 109.270 318.750 109.560 ;
        RECT 320.800 109.220 322.000 109.510 ;
        RECT 323.510 109.190 326.135 109.600 ;
        RECT 327.720 109.285 328.100 109.665 ;
        RECT 363.805 109.595 367.065 109.975 ;
        RECT 367.805 109.595 371.065 109.975 ;
        RECT 377.305 109.595 380.565 109.975 ;
        RECT 381.305 109.595 384.565 109.975 ;
        RECT 314.755 108.510 330.675 108.810 ;
        RECT 315.290 107.765 332.235 108.065 ;
        RECT 364.470 107.680 390.765 108.020 ;
        RECT 325.695 106.750 333.395 107.025 ;
        RECT 396.900 106.920 397.280 114.080 ;
        RECT 398.730 109.865 402.105 110.265 ;
        RECT 402.475 109.625 402.855 110.005 ;
        RECT 405.190 109.665 405.570 110.045 ;
        RECT 409.375 109.615 409.755 109.995 ;
        RECT 399.800 109.200 401.540 109.490 ;
        RECT 403.590 109.150 404.790 109.440 ;
        RECT 406.300 109.120 408.910 109.545 ;
        RECT 410.510 109.215 410.890 109.595 ;
        RECT 398.045 108.440 411.610 108.755 ;
        RECT 398.040 107.695 411.600 107.995 ;
        RECT 398.060 106.980 404.785 107.280 ;
        RECT 408.485 106.680 411.590 106.955 ;
        RECT 412.360 106.920 412.740 114.080 ;
        RECT 465.800 113.095 494.575 113.115 ;
        RECT 429.000 112.830 494.575 113.095 ;
        RECT 429.000 112.810 466.550 112.830 ;
        RECT 496.245 112.810 502.950 113.110 ;
        RECT 430.510 111.900 431.965 112.280 ;
        RECT 432.705 111.900 433.905 112.280 ;
        RECT 435.660 111.685 437.935 112.195 ;
        RECT 440.560 111.685 442.860 112.195 ;
        RECT 445.155 111.685 447.435 112.195 ;
        RECT 452.230 112.000 453.465 112.380 ;
        RECT 454.205 112.000 455.485 112.380 ;
        RECT 469.105 111.920 470.560 112.300 ;
        RECT 474.255 111.705 476.530 112.215 ;
        RECT 479.155 111.705 481.455 112.215 ;
        RECT 483.750 111.705 486.030 112.215 ;
        RECT 492.800 112.020 494.080 112.400 ;
        RECT 453.645 111.645 454.025 111.680 ;
        RECT 492.240 111.665 492.620 111.700 ;
        RECT 432.145 111.540 432.525 111.580 ;
        RECT 432.075 111.235 434.910 111.540 ;
        RECT 450.890 111.335 454.025 111.645 ;
        RECT 470.740 111.560 471.120 111.600 ;
        RECT 453.645 111.300 454.025 111.335 ;
        RECT 470.670 111.255 473.505 111.560 ;
        RECT 489.485 111.355 492.620 111.665 ;
        RECT 492.240 111.320 492.620 111.355 ;
        RECT 432.145 111.200 432.525 111.235 ;
        RECT 470.740 111.220 471.120 111.255 ;
        RECT 414.190 109.825 417.595 110.265 ;
        RECT 417.935 109.625 418.315 110.005 ;
        RECT 420.650 109.665 421.030 110.045 ;
        RECT 424.835 109.615 425.215 109.995 ;
        RECT 430.670 109.600 431.965 109.980 ;
        RECT 432.705 109.600 435.965 109.980 ;
        RECT 436.705 109.600 439.965 109.980 ;
        RECT 440.705 109.600 441.890 109.980 ;
        RECT 444.155 109.600 445.465 109.980 ;
        RECT 446.205 109.600 449.465 109.980 ;
        RECT 450.205 109.600 453.465 109.980 ;
        RECT 454.205 109.600 455.220 109.980 ;
        RECT 469.265 109.620 470.560 110.000 ;
        RECT 475.300 109.620 478.560 110.000 ;
        RECT 479.300 109.620 480.485 110.000 ;
        RECT 482.750 109.620 484.060 110.000 ;
        RECT 484.800 109.620 488.060 110.000 ;
        RECT 492.800 109.620 493.815 110.000 ;
        RECT 496.880 109.865 500.295 110.285 ;
        RECT 500.625 109.645 501.005 110.025 ;
        RECT 503.340 109.685 503.720 110.065 ;
        RECT 507.525 109.635 507.905 110.015 ;
        RECT 415.260 109.200 417.000 109.490 ;
        RECT 419.050 109.150 420.250 109.440 ;
        RECT 421.760 109.120 424.355 109.495 ;
        RECT 425.970 109.215 426.350 109.595 ;
        RECT 432.145 108.900 432.525 109.280 ;
        RECT 436.145 108.900 436.525 109.280 ;
        RECT 440.145 109.235 440.525 109.280 ;
        RECT 445.645 109.235 446.025 109.280 ;
        RECT 440.095 108.920 446.030 109.235 ;
        RECT 440.145 108.900 440.525 108.920 ;
        RECT 445.645 108.900 446.025 108.920 ;
        RECT 449.645 108.900 450.025 109.280 ;
        RECT 453.645 108.900 454.025 109.280 ;
        RECT 470.740 108.920 471.120 109.300 ;
        RECT 474.740 108.920 475.120 109.300 ;
        RECT 478.740 109.255 479.120 109.300 ;
        RECT 484.240 109.255 484.620 109.300 ;
        RECT 478.690 108.940 484.625 109.255 ;
        RECT 478.740 108.920 479.120 108.940 ;
        RECT 484.240 108.920 484.620 108.940 ;
        RECT 488.240 108.920 488.620 109.300 ;
        RECT 492.240 108.920 492.620 109.300 ;
        RECT 497.950 109.220 499.690 109.510 ;
        RECT 501.740 109.170 502.940 109.460 ;
        RECT 504.450 109.130 507.080 109.585 ;
        RECT 508.660 109.235 509.040 109.615 ;
        RECT 413.500 108.440 427.325 108.740 ;
        RECT 429.000 108.275 445.010 108.650 ;
        RECT 462.830 108.295 483.605 108.670 ;
        RECT 413.505 107.695 431.925 107.995 ;
        RECT 433.370 107.685 460.680 108.025 ;
        RECT 412.985 106.980 420.245 107.280 ;
        RECT 262.305 106.625 289.865 106.635 ;
        RECT 232.600 106.605 251.270 106.615 ;
        RECT 262.305 106.605 298.870 106.625 ;
        RECT 232.600 106.315 298.870 106.605 ;
        RECT 398.040 106.360 402.165 106.630 ;
        RECT 413.540 106.445 417.625 106.715 ;
        RECT 423.945 106.680 427.695 106.955 ;
        RECT 429.000 106.920 455.230 107.310 ;
        RECT 461.860 106.940 493.825 107.330 ;
        RECT 506.635 106.700 509.765 106.975 ;
        RECT 510.510 106.940 510.890 114.100 ;
        RECT 560.125 111.940 561.325 112.320 ;
        RECT 511.750 111.640 518.490 111.940 ;
        RECT 563.080 111.725 565.355 112.235 ;
        RECT 567.980 111.725 570.280 112.235 ;
        RECT 572.575 111.725 574.855 112.235 ;
        RECT 579.650 112.040 580.885 112.420 ;
        RECT 512.340 109.845 515.795 110.285 ;
        RECT 516.085 109.645 516.465 110.025 ;
        RECT 518.800 109.685 519.180 110.065 ;
        RECT 522.985 109.635 523.365 110.015 ;
        RECT 560.125 109.640 563.385 110.020 ;
        RECT 564.125 109.640 567.385 110.020 ;
        RECT 573.625 109.640 576.885 110.020 ;
        RECT 577.625 109.640 580.885 110.020 ;
        RECT 513.410 109.220 515.150 109.510 ;
        RECT 517.200 109.170 518.400 109.460 ;
        RECT 519.910 109.140 522.535 109.550 ;
        RECT 524.120 109.235 524.500 109.615 ;
        RECT 511.155 108.460 527.075 108.760 ;
        RECT 511.690 107.715 528.635 108.015 ;
        RECT 560.790 107.725 587.085 108.065 ;
        RECT 522.095 106.700 529.795 106.975 ;
        RECT 593.275 106.955 593.655 114.115 ;
        RECT 595.105 109.900 598.480 110.300 ;
        RECT 598.850 109.660 599.230 110.040 ;
        RECT 601.565 109.700 601.945 110.080 ;
        RECT 605.750 109.650 606.130 110.030 ;
        RECT 596.175 109.235 597.915 109.525 ;
        RECT 599.965 109.185 601.165 109.475 ;
        RECT 602.675 109.155 605.285 109.580 ;
        RECT 606.885 109.250 607.265 109.630 ;
        RECT 594.420 108.475 607.985 108.790 ;
        RECT 594.415 107.730 607.975 108.030 ;
        RECT 594.435 107.015 601.160 107.315 ;
        RECT 604.860 106.715 607.965 106.990 ;
        RECT 608.735 106.955 609.115 114.115 ;
        RECT 662.175 113.130 690.950 113.150 ;
        RECT 625.375 112.865 690.950 113.130 ;
        RECT 625.375 112.845 662.925 112.865 ;
        RECT 692.620 112.845 699.325 113.145 ;
        RECT 626.885 111.935 628.340 112.315 ;
        RECT 629.080 111.935 630.280 112.315 ;
        RECT 632.035 111.720 634.310 112.230 ;
        RECT 636.935 111.720 639.235 112.230 ;
        RECT 641.530 111.720 643.810 112.230 ;
        RECT 648.605 112.035 649.840 112.415 ;
        RECT 650.580 112.035 651.860 112.415 ;
        RECT 665.480 111.955 666.935 112.335 ;
        RECT 670.630 111.740 672.905 112.250 ;
        RECT 675.530 111.740 677.830 112.250 ;
        RECT 680.125 111.740 682.405 112.250 ;
        RECT 689.175 112.055 690.455 112.435 ;
        RECT 650.020 111.680 650.400 111.715 ;
        RECT 688.615 111.700 688.995 111.735 ;
        RECT 628.520 111.575 628.900 111.615 ;
        RECT 628.450 111.270 631.285 111.575 ;
        RECT 647.265 111.370 650.400 111.680 ;
        RECT 667.115 111.595 667.495 111.635 ;
        RECT 650.020 111.335 650.400 111.370 ;
        RECT 667.045 111.290 669.880 111.595 ;
        RECT 685.860 111.390 688.995 111.700 ;
        RECT 688.615 111.355 688.995 111.390 ;
        RECT 628.520 111.235 628.900 111.270 ;
        RECT 667.115 111.255 667.495 111.290 ;
        RECT 610.565 109.860 613.970 110.300 ;
        RECT 614.310 109.660 614.690 110.040 ;
        RECT 617.025 109.700 617.405 110.080 ;
        RECT 621.210 109.650 621.590 110.030 ;
        RECT 627.045 109.635 628.340 110.015 ;
        RECT 629.080 109.635 632.340 110.015 ;
        RECT 633.080 109.635 636.340 110.015 ;
        RECT 637.080 109.635 638.265 110.015 ;
        RECT 640.530 109.635 641.840 110.015 ;
        RECT 642.580 109.635 645.840 110.015 ;
        RECT 646.580 109.635 649.840 110.015 ;
        RECT 650.580 109.635 651.595 110.015 ;
        RECT 665.640 109.655 666.935 110.035 ;
        RECT 671.675 109.655 674.935 110.035 ;
        RECT 675.675 109.655 676.860 110.035 ;
        RECT 679.125 109.655 680.435 110.035 ;
        RECT 681.175 109.655 684.435 110.035 ;
        RECT 689.175 109.655 690.190 110.035 ;
        RECT 693.255 109.900 696.670 110.320 ;
        RECT 697.000 109.680 697.380 110.060 ;
        RECT 699.715 109.720 700.095 110.100 ;
        RECT 703.900 109.670 704.280 110.050 ;
        RECT 611.635 109.235 613.375 109.525 ;
        RECT 615.425 109.185 616.625 109.475 ;
        RECT 618.135 109.155 620.730 109.530 ;
        RECT 622.345 109.250 622.725 109.630 ;
        RECT 628.520 108.935 628.900 109.315 ;
        RECT 632.520 108.935 632.900 109.315 ;
        RECT 636.520 109.270 636.900 109.315 ;
        RECT 642.020 109.270 642.400 109.315 ;
        RECT 636.470 108.955 642.405 109.270 ;
        RECT 636.520 108.935 636.900 108.955 ;
        RECT 642.020 108.935 642.400 108.955 ;
        RECT 646.020 108.935 646.400 109.315 ;
        RECT 650.020 108.935 650.400 109.315 ;
        RECT 667.115 108.955 667.495 109.335 ;
        RECT 671.115 108.955 671.495 109.335 ;
        RECT 675.115 109.290 675.495 109.335 ;
        RECT 680.615 109.290 680.995 109.335 ;
        RECT 675.065 108.975 681.000 109.290 ;
        RECT 675.115 108.955 675.495 108.975 ;
        RECT 680.615 108.955 680.995 108.975 ;
        RECT 684.615 108.955 684.995 109.335 ;
        RECT 688.615 108.955 688.995 109.335 ;
        RECT 694.325 109.255 696.065 109.545 ;
        RECT 698.115 109.205 699.315 109.495 ;
        RECT 700.825 109.165 703.455 109.620 ;
        RECT 705.035 109.270 705.415 109.650 ;
        RECT 609.875 108.475 623.700 108.775 ;
        RECT 625.375 108.310 641.385 108.685 ;
        RECT 659.205 108.330 679.980 108.705 ;
        RECT 609.880 107.730 628.300 108.030 ;
        RECT 629.745 107.720 657.055 108.060 ;
        RECT 609.360 107.015 616.620 107.315 ;
        RECT 458.705 106.575 486.265 106.585 ;
        RECT 429.000 106.555 447.670 106.565 ;
        RECT 458.705 106.555 495.270 106.575 ;
        RECT 36.235 106.295 66.255 106.315 ;
        RECT 232.600 106.295 262.620 106.315 ;
        RECT 429.000 106.265 495.270 106.555 ;
        RECT 594.415 106.395 598.540 106.665 ;
        RECT 609.915 106.480 614.000 106.750 ;
        RECT 620.320 106.715 624.070 106.990 ;
        RECT 625.375 106.955 651.605 107.345 ;
        RECT 658.235 106.975 690.200 107.365 ;
        RECT 703.010 106.735 706.140 107.010 ;
        RECT 706.885 106.975 707.265 114.135 ;
        RECT 754.005 114.125 779.440 115.025 ;
        RECT 861.530 115.015 917.885 115.035 ;
        RECT 1057.870 115.015 1114.225 115.035 ;
        RECT 1254.210 115.015 1310.565 115.035 ;
        RECT 789.245 114.135 917.885 115.015 ;
        RECT 789.245 114.115 861.635 114.135 ;
        RECT 708.125 111.675 714.865 111.975 ;
        RECT 756.490 111.945 757.690 112.325 ;
        RECT 759.445 111.730 761.720 112.240 ;
        RECT 764.345 111.730 766.645 112.240 ;
        RECT 768.940 111.730 771.220 112.240 ;
        RECT 776.015 112.045 777.250 112.425 ;
        RECT 708.715 109.880 712.170 110.320 ;
        RECT 712.460 109.680 712.840 110.060 ;
        RECT 715.175 109.720 715.555 110.100 ;
        RECT 719.360 109.670 719.740 110.050 ;
        RECT 709.785 109.255 711.525 109.545 ;
        RECT 713.575 109.205 714.775 109.495 ;
        RECT 716.285 109.175 718.910 109.585 ;
        RECT 720.495 109.270 720.875 109.650 ;
        RECT 756.490 109.645 759.750 110.025 ;
        RECT 760.490 109.645 763.750 110.025 ;
        RECT 769.990 109.645 773.250 110.025 ;
        RECT 773.990 109.645 777.250 110.025 ;
        RECT 707.530 108.495 723.450 108.795 ;
        RECT 708.065 107.750 725.010 108.050 ;
        RECT 757.155 107.730 783.450 108.070 ;
        RECT 718.470 106.735 726.170 107.010 ;
        RECT 789.615 106.955 789.995 114.115 ;
        RECT 791.445 109.900 794.820 110.300 ;
        RECT 795.190 109.660 795.570 110.040 ;
        RECT 797.905 109.700 798.285 110.080 ;
        RECT 802.090 109.650 802.470 110.030 ;
        RECT 792.515 109.235 794.255 109.525 ;
        RECT 796.305 109.185 797.505 109.475 ;
        RECT 799.015 109.155 801.625 109.580 ;
        RECT 803.225 109.250 803.605 109.630 ;
        RECT 790.760 108.475 804.325 108.790 ;
        RECT 790.755 107.730 804.315 108.030 ;
        RECT 790.775 107.015 797.500 107.315 ;
        RECT 801.200 106.715 804.305 106.990 ;
        RECT 805.075 106.955 805.455 114.115 ;
        RECT 858.515 113.130 887.290 113.150 ;
        RECT 821.715 112.865 887.290 113.130 ;
        RECT 821.715 112.845 859.265 112.865 ;
        RECT 888.960 112.845 895.665 113.145 ;
        RECT 823.225 111.935 824.680 112.315 ;
        RECT 825.420 111.935 826.620 112.315 ;
        RECT 828.375 111.720 830.650 112.230 ;
        RECT 833.275 111.720 835.575 112.230 ;
        RECT 837.870 111.720 840.150 112.230 ;
        RECT 844.945 112.035 846.180 112.415 ;
        RECT 846.920 112.035 848.200 112.415 ;
        RECT 861.820 111.955 863.275 112.335 ;
        RECT 866.970 111.740 869.245 112.250 ;
        RECT 871.870 111.740 874.170 112.250 ;
        RECT 876.465 111.740 878.745 112.250 ;
        RECT 885.515 112.055 886.795 112.435 ;
        RECT 846.360 111.680 846.740 111.715 ;
        RECT 884.955 111.700 885.335 111.735 ;
        RECT 824.860 111.575 825.240 111.615 ;
        RECT 824.790 111.270 827.625 111.575 ;
        RECT 843.605 111.370 846.740 111.680 ;
        RECT 863.455 111.595 863.835 111.635 ;
        RECT 846.360 111.335 846.740 111.370 ;
        RECT 863.385 111.290 866.220 111.595 ;
        RECT 882.200 111.390 885.335 111.700 ;
        RECT 884.955 111.355 885.335 111.390 ;
        RECT 824.860 111.235 825.240 111.270 ;
        RECT 863.455 111.255 863.835 111.290 ;
        RECT 806.905 109.860 810.310 110.300 ;
        RECT 810.650 109.660 811.030 110.040 ;
        RECT 813.365 109.700 813.745 110.080 ;
        RECT 817.550 109.650 817.930 110.030 ;
        RECT 823.385 109.635 824.680 110.015 ;
        RECT 825.420 109.635 828.680 110.015 ;
        RECT 829.420 109.635 832.680 110.015 ;
        RECT 833.420 109.635 834.605 110.015 ;
        RECT 836.870 109.635 838.180 110.015 ;
        RECT 838.920 109.635 842.180 110.015 ;
        RECT 842.920 109.635 846.180 110.015 ;
        RECT 846.920 109.635 847.935 110.015 ;
        RECT 861.980 109.655 863.275 110.035 ;
        RECT 868.015 109.655 871.275 110.035 ;
        RECT 872.015 109.655 873.200 110.035 ;
        RECT 875.465 109.655 876.775 110.035 ;
        RECT 877.515 109.655 880.775 110.035 ;
        RECT 885.515 109.655 886.530 110.035 ;
        RECT 889.595 109.900 893.010 110.320 ;
        RECT 893.340 109.680 893.720 110.060 ;
        RECT 896.055 109.720 896.435 110.100 ;
        RECT 900.240 109.670 900.620 110.050 ;
        RECT 807.975 109.235 809.715 109.525 ;
        RECT 811.765 109.185 812.965 109.475 ;
        RECT 814.475 109.155 817.070 109.530 ;
        RECT 818.685 109.250 819.065 109.630 ;
        RECT 824.860 108.935 825.240 109.315 ;
        RECT 828.860 108.935 829.240 109.315 ;
        RECT 832.860 109.270 833.240 109.315 ;
        RECT 838.360 109.270 838.740 109.315 ;
        RECT 832.810 108.955 838.745 109.270 ;
        RECT 832.860 108.935 833.240 108.955 ;
        RECT 838.360 108.935 838.740 108.955 ;
        RECT 842.360 108.935 842.740 109.315 ;
        RECT 846.360 108.935 846.740 109.315 ;
        RECT 863.455 108.955 863.835 109.335 ;
        RECT 867.455 108.955 867.835 109.335 ;
        RECT 871.455 109.290 871.835 109.335 ;
        RECT 876.955 109.290 877.335 109.335 ;
        RECT 871.405 108.975 877.340 109.290 ;
        RECT 871.455 108.955 871.835 108.975 ;
        RECT 876.955 108.955 877.335 108.975 ;
        RECT 880.955 108.955 881.335 109.335 ;
        RECT 884.955 108.955 885.335 109.335 ;
        RECT 890.665 109.255 892.405 109.545 ;
        RECT 894.455 109.205 895.655 109.495 ;
        RECT 897.165 109.165 899.795 109.620 ;
        RECT 901.375 109.270 901.755 109.650 ;
        RECT 806.215 108.475 820.040 108.775 ;
        RECT 821.715 108.310 837.725 108.685 ;
        RECT 855.545 108.330 876.320 108.705 ;
        RECT 806.220 107.730 824.640 108.030 ;
        RECT 826.085 107.720 853.395 108.060 ;
        RECT 805.700 107.015 812.960 107.315 ;
        RECT 655.080 106.610 682.640 106.620 ;
        RECT 625.375 106.590 644.045 106.600 ;
        RECT 655.080 106.590 691.645 106.610 ;
        RECT 625.375 106.300 691.645 106.590 ;
        RECT 790.755 106.395 794.880 106.665 ;
        RECT 806.255 106.480 810.340 106.750 ;
        RECT 816.660 106.715 820.410 106.990 ;
        RECT 821.715 106.955 847.945 107.345 ;
        RECT 854.575 106.975 886.540 107.365 ;
        RECT 899.350 106.735 902.480 107.010 ;
        RECT 903.225 106.975 903.605 114.135 ;
        RECT 950.390 114.110 975.825 115.010 ;
        RECT 985.585 114.135 1114.225 115.015 ;
        RECT 985.585 114.115 1057.975 114.135 ;
        RECT 904.465 111.675 911.205 111.975 ;
        RECT 952.875 111.930 954.075 112.310 ;
        RECT 955.830 111.715 958.105 112.225 ;
        RECT 960.730 111.715 963.030 112.225 ;
        RECT 965.325 111.715 967.605 112.225 ;
        RECT 972.400 112.030 973.635 112.410 ;
        RECT 905.055 109.880 908.510 110.320 ;
        RECT 908.800 109.680 909.180 110.060 ;
        RECT 911.515 109.720 911.895 110.100 ;
        RECT 915.700 109.670 916.080 110.050 ;
        RECT 906.125 109.255 907.865 109.545 ;
        RECT 909.915 109.205 911.115 109.495 ;
        RECT 912.625 109.175 915.250 109.585 ;
        RECT 916.835 109.270 917.215 109.650 ;
        RECT 952.875 109.630 956.135 110.010 ;
        RECT 956.875 109.630 960.135 110.010 ;
        RECT 966.375 109.630 969.635 110.010 ;
        RECT 970.375 109.630 973.635 110.010 ;
        RECT 903.870 108.495 919.790 108.795 ;
        RECT 904.405 107.750 921.350 108.050 ;
        RECT 953.540 107.715 979.835 108.055 ;
        RECT 914.810 106.735 922.510 107.010 ;
        RECT 985.955 106.955 986.335 114.115 ;
        RECT 987.785 109.900 991.160 110.300 ;
        RECT 991.530 109.660 991.910 110.040 ;
        RECT 994.245 109.700 994.625 110.080 ;
        RECT 998.430 109.650 998.810 110.030 ;
        RECT 988.855 109.235 990.595 109.525 ;
        RECT 992.645 109.185 993.845 109.475 ;
        RECT 995.355 109.155 997.965 109.580 ;
        RECT 999.565 109.250 999.945 109.630 ;
        RECT 987.100 108.475 1000.665 108.790 ;
        RECT 987.095 107.730 1000.655 108.030 ;
        RECT 987.115 107.015 993.840 107.315 ;
        RECT 997.540 106.715 1000.645 106.990 ;
        RECT 1001.415 106.955 1001.795 114.115 ;
        RECT 1054.855 113.130 1083.630 113.150 ;
        RECT 1018.055 112.865 1083.630 113.130 ;
        RECT 1018.055 112.845 1055.605 112.865 ;
        RECT 1085.300 112.845 1092.005 113.145 ;
        RECT 1019.565 111.935 1021.020 112.315 ;
        RECT 1021.760 111.935 1022.960 112.315 ;
        RECT 1024.715 111.720 1026.990 112.230 ;
        RECT 1029.615 111.720 1031.915 112.230 ;
        RECT 1034.210 111.720 1036.490 112.230 ;
        RECT 1041.285 112.035 1042.520 112.415 ;
        RECT 1043.260 112.035 1044.540 112.415 ;
        RECT 1058.160 111.955 1059.615 112.335 ;
        RECT 1063.310 111.740 1065.585 112.250 ;
        RECT 1068.210 111.740 1070.510 112.250 ;
        RECT 1072.805 111.740 1075.085 112.250 ;
        RECT 1081.855 112.055 1083.135 112.435 ;
        RECT 1042.700 111.680 1043.080 111.715 ;
        RECT 1081.295 111.700 1081.675 111.735 ;
        RECT 1021.200 111.575 1021.580 111.615 ;
        RECT 1021.130 111.270 1023.965 111.575 ;
        RECT 1039.945 111.370 1043.080 111.680 ;
        RECT 1059.795 111.595 1060.175 111.635 ;
        RECT 1042.700 111.335 1043.080 111.370 ;
        RECT 1059.725 111.290 1062.560 111.595 ;
        RECT 1078.540 111.390 1081.675 111.700 ;
        RECT 1081.295 111.355 1081.675 111.390 ;
        RECT 1021.200 111.235 1021.580 111.270 ;
        RECT 1059.795 111.255 1060.175 111.290 ;
        RECT 1003.245 109.860 1006.650 110.300 ;
        RECT 1006.990 109.660 1007.370 110.040 ;
        RECT 1009.705 109.700 1010.085 110.080 ;
        RECT 1013.890 109.650 1014.270 110.030 ;
        RECT 1019.725 109.635 1021.020 110.015 ;
        RECT 1021.760 109.635 1025.020 110.015 ;
        RECT 1025.760 109.635 1029.020 110.015 ;
        RECT 1029.760 109.635 1030.945 110.015 ;
        RECT 1033.210 109.635 1034.520 110.015 ;
        RECT 1035.260 109.635 1038.520 110.015 ;
        RECT 1039.260 109.635 1042.520 110.015 ;
        RECT 1043.260 109.635 1044.275 110.015 ;
        RECT 1058.320 109.655 1059.615 110.035 ;
        RECT 1064.355 109.655 1067.615 110.035 ;
        RECT 1068.355 109.655 1069.540 110.035 ;
        RECT 1071.805 109.655 1073.115 110.035 ;
        RECT 1073.855 109.655 1077.115 110.035 ;
        RECT 1081.855 109.655 1082.870 110.035 ;
        RECT 1085.935 109.900 1089.350 110.320 ;
        RECT 1089.680 109.680 1090.060 110.060 ;
        RECT 1092.395 109.720 1092.775 110.100 ;
        RECT 1096.580 109.670 1096.960 110.050 ;
        RECT 1004.315 109.235 1006.055 109.525 ;
        RECT 1008.105 109.185 1009.305 109.475 ;
        RECT 1010.815 109.155 1013.410 109.530 ;
        RECT 1015.025 109.250 1015.405 109.630 ;
        RECT 1021.200 108.935 1021.580 109.315 ;
        RECT 1025.200 108.935 1025.580 109.315 ;
        RECT 1029.200 109.270 1029.580 109.315 ;
        RECT 1034.700 109.270 1035.080 109.315 ;
        RECT 1029.150 108.955 1035.085 109.270 ;
        RECT 1029.200 108.935 1029.580 108.955 ;
        RECT 1034.700 108.935 1035.080 108.955 ;
        RECT 1038.700 108.935 1039.080 109.315 ;
        RECT 1042.700 108.935 1043.080 109.315 ;
        RECT 1059.795 108.955 1060.175 109.335 ;
        RECT 1063.795 108.955 1064.175 109.335 ;
        RECT 1067.795 109.290 1068.175 109.335 ;
        RECT 1073.295 109.290 1073.675 109.335 ;
        RECT 1067.745 108.975 1073.680 109.290 ;
        RECT 1067.795 108.955 1068.175 108.975 ;
        RECT 1073.295 108.955 1073.675 108.975 ;
        RECT 1077.295 108.955 1077.675 109.335 ;
        RECT 1081.295 108.955 1081.675 109.335 ;
        RECT 1087.005 109.255 1088.745 109.545 ;
        RECT 1090.795 109.205 1091.995 109.495 ;
        RECT 1093.505 109.165 1096.135 109.620 ;
        RECT 1097.715 109.270 1098.095 109.650 ;
        RECT 1002.555 108.475 1016.380 108.775 ;
        RECT 1018.055 108.310 1034.065 108.685 ;
        RECT 1051.885 108.330 1072.660 108.705 ;
        RECT 1002.560 107.730 1020.980 108.030 ;
        RECT 1022.425 107.720 1049.735 108.060 ;
        RECT 1002.040 107.015 1009.300 107.315 ;
        RECT 851.420 106.610 878.980 106.620 ;
        RECT 821.715 106.590 840.385 106.600 ;
        RECT 851.420 106.590 887.985 106.610 ;
        RECT 821.715 106.300 887.985 106.590 ;
        RECT 987.095 106.395 991.220 106.665 ;
        RECT 1002.595 106.480 1006.680 106.750 ;
        RECT 1013.000 106.715 1016.750 106.990 ;
        RECT 1018.055 106.955 1044.285 107.345 ;
        RECT 1050.915 106.975 1082.880 107.365 ;
        RECT 1095.690 106.735 1098.820 107.010 ;
        RECT 1099.565 106.975 1099.945 114.135 ;
        RECT 1146.715 114.115 1172.150 115.015 ;
        RECT 1181.925 114.135 1310.565 115.015 ;
        RECT 1181.925 114.115 1254.315 114.135 ;
        RECT 1100.805 111.675 1107.545 111.975 ;
        RECT 1149.200 111.935 1150.400 112.315 ;
        RECT 1152.155 111.720 1154.430 112.230 ;
        RECT 1157.055 111.720 1159.355 112.230 ;
        RECT 1161.650 111.720 1163.930 112.230 ;
        RECT 1168.725 112.035 1169.960 112.415 ;
        RECT 1101.395 109.880 1104.850 110.320 ;
        RECT 1105.140 109.680 1105.520 110.060 ;
        RECT 1107.855 109.720 1108.235 110.100 ;
        RECT 1112.040 109.670 1112.420 110.050 ;
        RECT 1102.465 109.255 1104.205 109.545 ;
        RECT 1106.255 109.205 1107.455 109.495 ;
        RECT 1108.965 109.175 1111.590 109.585 ;
        RECT 1113.175 109.270 1113.555 109.650 ;
        RECT 1149.200 109.635 1152.460 110.015 ;
        RECT 1153.200 109.635 1156.460 110.015 ;
        RECT 1162.700 109.635 1165.960 110.015 ;
        RECT 1166.700 109.635 1169.960 110.015 ;
        RECT 1100.210 108.495 1116.130 108.795 ;
        RECT 1100.745 107.750 1117.690 108.050 ;
        RECT 1149.865 107.720 1176.160 108.060 ;
        RECT 1111.150 106.735 1118.850 107.010 ;
        RECT 1182.295 106.955 1182.675 114.115 ;
        RECT 1184.125 109.900 1187.500 110.300 ;
        RECT 1187.870 109.660 1188.250 110.040 ;
        RECT 1190.585 109.700 1190.965 110.080 ;
        RECT 1194.770 109.650 1195.150 110.030 ;
        RECT 1185.195 109.235 1186.935 109.525 ;
        RECT 1188.985 109.185 1190.185 109.475 ;
        RECT 1191.695 109.155 1194.305 109.580 ;
        RECT 1195.905 109.250 1196.285 109.630 ;
        RECT 1183.440 108.475 1197.005 108.790 ;
        RECT 1183.435 107.730 1196.995 108.030 ;
        RECT 1183.455 107.015 1190.180 107.315 ;
        RECT 1193.880 106.715 1196.985 106.990 ;
        RECT 1197.755 106.955 1198.135 114.115 ;
        RECT 1251.195 113.130 1279.970 113.150 ;
        RECT 1214.395 112.865 1279.970 113.130 ;
        RECT 1214.395 112.845 1251.945 112.865 ;
        RECT 1281.640 112.845 1288.345 113.145 ;
        RECT 1215.905 111.935 1217.360 112.315 ;
        RECT 1218.100 111.935 1219.300 112.315 ;
        RECT 1221.055 111.720 1223.330 112.230 ;
        RECT 1225.955 111.720 1228.255 112.230 ;
        RECT 1230.550 111.720 1232.830 112.230 ;
        RECT 1237.625 112.035 1238.860 112.415 ;
        RECT 1239.600 112.035 1240.880 112.415 ;
        RECT 1254.500 111.955 1255.955 112.335 ;
        RECT 1256.695 111.955 1257.895 112.335 ;
        RECT 1259.650 111.740 1261.925 112.250 ;
        RECT 1264.550 111.740 1266.850 112.250 ;
        RECT 1269.145 111.740 1271.425 112.250 ;
        RECT 1276.220 112.055 1277.455 112.435 ;
        RECT 1278.195 112.055 1279.475 112.435 ;
        RECT 1239.040 111.680 1239.420 111.715 ;
        RECT 1277.635 111.700 1278.015 111.735 ;
        RECT 1217.540 111.575 1217.920 111.615 ;
        RECT 1217.470 111.270 1220.305 111.575 ;
        RECT 1236.285 111.370 1239.420 111.680 ;
        RECT 1256.135 111.595 1256.515 111.635 ;
        RECT 1239.040 111.335 1239.420 111.370 ;
        RECT 1256.065 111.290 1258.900 111.595 ;
        RECT 1274.880 111.390 1278.015 111.700 ;
        RECT 1277.635 111.355 1278.015 111.390 ;
        RECT 1217.540 111.235 1217.920 111.270 ;
        RECT 1256.135 111.255 1256.515 111.290 ;
        RECT 1199.585 109.860 1202.990 110.300 ;
        RECT 1203.330 109.660 1203.710 110.040 ;
        RECT 1206.045 109.700 1206.425 110.080 ;
        RECT 1210.230 109.650 1210.610 110.030 ;
        RECT 1216.065 109.635 1217.360 110.015 ;
        RECT 1218.100 109.635 1221.360 110.015 ;
        RECT 1222.100 109.635 1225.360 110.015 ;
        RECT 1226.100 109.635 1227.285 110.015 ;
        RECT 1229.550 109.635 1230.860 110.015 ;
        RECT 1231.600 109.635 1234.860 110.015 ;
        RECT 1235.600 109.635 1238.860 110.015 ;
        RECT 1239.600 109.635 1240.615 110.015 ;
        RECT 1254.660 109.655 1255.955 110.035 ;
        RECT 1256.695 109.655 1259.955 110.035 ;
        RECT 1260.695 109.655 1263.955 110.035 ;
        RECT 1264.695 109.655 1265.880 110.035 ;
        RECT 1268.145 109.655 1269.455 110.035 ;
        RECT 1270.195 109.655 1273.455 110.035 ;
        RECT 1274.195 109.655 1277.455 110.035 ;
        RECT 1278.195 109.655 1279.210 110.035 ;
        RECT 1282.275 109.900 1285.690 110.320 ;
        RECT 1286.020 109.680 1286.400 110.060 ;
        RECT 1288.735 109.720 1289.115 110.100 ;
        RECT 1292.920 109.670 1293.300 110.050 ;
        RECT 1200.655 109.235 1202.395 109.525 ;
        RECT 1204.445 109.185 1205.645 109.475 ;
        RECT 1207.155 109.155 1209.750 109.530 ;
        RECT 1211.365 109.250 1211.745 109.630 ;
        RECT 1217.540 108.935 1217.920 109.315 ;
        RECT 1221.540 108.935 1221.920 109.315 ;
        RECT 1225.540 109.270 1225.920 109.315 ;
        RECT 1231.040 109.270 1231.420 109.315 ;
        RECT 1225.490 108.955 1231.425 109.270 ;
        RECT 1225.540 108.935 1225.920 108.955 ;
        RECT 1231.040 108.935 1231.420 108.955 ;
        RECT 1235.040 108.935 1235.420 109.315 ;
        RECT 1239.040 108.935 1239.420 109.315 ;
        RECT 1256.135 108.955 1256.515 109.335 ;
        RECT 1260.135 108.955 1260.515 109.335 ;
        RECT 1264.135 109.290 1264.515 109.335 ;
        RECT 1269.635 109.290 1270.015 109.335 ;
        RECT 1264.085 108.975 1270.020 109.290 ;
        RECT 1264.135 108.955 1264.515 108.975 ;
        RECT 1269.635 108.955 1270.015 108.975 ;
        RECT 1273.635 108.955 1274.015 109.335 ;
        RECT 1277.635 108.955 1278.015 109.335 ;
        RECT 1283.345 109.255 1285.085 109.545 ;
        RECT 1287.135 109.205 1288.335 109.495 ;
        RECT 1289.845 109.165 1292.475 109.620 ;
        RECT 1294.055 109.270 1294.435 109.650 ;
        RECT 1198.895 108.475 1212.720 108.775 ;
        RECT 1214.395 108.310 1230.405 108.685 ;
        RECT 1248.225 108.330 1269.000 108.705 ;
        RECT 1281.625 108.495 1295.240 108.795 ;
        RECT 1198.900 107.730 1217.320 108.030 ;
        RECT 1218.765 107.720 1246.075 108.060 ;
        RECT 1257.360 107.740 1279.915 108.080 ;
        RECT 1281.025 107.750 1295.670 108.050 ;
        RECT 1198.380 107.015 1205.640 107.315 ;
        RECT 1047.760 106.610 1075.320 106.620 ;
        RECT 1018.055 106.590 1036.725 106.600 ;
        RECT 1047.760 106.590 1084.325 106.610 ;
        RECT 1018.055 106.300 1084.325 106.590 ;
        RECT 1183.435 106.395 1187.560 106.665 ;
        RECT 1198.935 106.480 1203.020 106.750 ;
        RECT 1209.340 106.715 1213.090 106.990 ;
        RECT 1214.395 106.955 1240.625 107.345 ;
        RECT 1247.255 106.975 1279.220 107.365 ;
        RECT 1292.030 106.735 1295.160 107.010 ;
        RECT 1295.905 106.975 1296.285 114.135 ;
        RECT 1297.145 111.675 1303.885 111.975 ;
        RECT 1297.735 109.880 1301.190 110.320 ;
        RECT 1304.195 109.720 1304.575 110.100 ;
        RECT 1302.595 109.205 1303.795 109.495 ;
        RECT 1309.515 109.270 1309.895 109.650 ;
        RECT 1296.550 108.495 1312.470 108.795 ;
        RECT 1297.085 107.750 1314.030 108.050 ;
        RECT 1244.100 106.610 1271.660 106.620 ;
        RECT 1214.395 106.590 1233.065 106.600 ;
        RECT 1244.100 106.590 1280.665 106.610 ;
        RECT 1214.395 106.300 1280.665 106.590 ;
        RECT 625.375 106.280 655.395 106.300 ;
        RECT 821.715 106.280 851.735 106.300 ;
        RECT 1018.055 106.280 1048.075 106.300 ;
        RECT 1214.395 106.280 1244.415 106.300 ;
        RECT 429.000 106.245 459.020 106.265 ;
        RECT 6.510 105.835 10.640 106.135 ;
        RECT -59.695 105.010 -56.130 105.020 ;
        RECT -59.695 104.685 -55.335 105.010 ;
        RECT -9.370 104.765 -3.455 105.100 ;
        RECT -6.100 104.745 -3.455 104.765 ;
        RECT -56.290 104.675 -55.335 104.685 ;
        RECT -79.100 104.045 -75.800 104.425 ;
        RECT -75.100 104.045 -71.800 104.425 ;
        RECT -65.600 104.045 -62.300 104.425 ;
        RECT -61.600 104.045 -58.300 104.425 ;
        RECT -28.775 104.125 -25.475 104.505 ;
        RECT -24.775 104.125 -21.475 104.505 ;
        RECT -15.275 104.125 -11.975 104.505 ;
        RECT -11.275 104.125 -7.975 104.505 ;
        RECT -79.100 102.045 -77.815 102.425 ;
        RECT -59.785 102.045 -58.300 102.425 ;
        RECT -28.775 102.125 -27.490 102.505 ;
        RECT -9.460 102.125 -7.975 102.505 ;
        RECT -77.595 101.365 -76.075 101.725 ;
        RECT -27.270 101.445 -25.750 101.805 ;
        RECT 4.135 100.005 4.515 105.835 ;
        RECT 13.015 105.785 17.515 106.095 ;
        RECT 21.970 105.835 26.100 106.135 ;
        RECT 8.975 105.235 15.365 105.525 ;
        RECT 8.390 104.655 19.045 104.990 ;
        RECT 7.740 104.070 10.660 104.370 ;
        RECT 14.205 104.055 17.575 104.355 ;
        RECT 5.955 103.320 6.335 103.700 ;
        RECT 8.360 103.335 10.140 103.625 ;
        RECT 11.615 103.425 12.805 103.710 ;
        RECT 15.735 103.305 17.045 103.625 ;
        RECT 7.090 102.720 7.470 103.100 ;
        RECT 10.835 102.760 11.215 103.140 ;
        RECT 13.545 102.750 13.925 103.130 ;
        RECT 14.955 102.595 18.135 102.915 ;
        RECT 4.885 100.005 8.980 100.010 ;
        RECT 19.595 100.005 19.975 105.835 ;
        RECT 28.475 105.785 32.975 106.095 ;
        RECT 120.120 105.855 124.250 106.155 ;
        RECT 71.160 105.625 102.905 105.645 ;
        RECT 24.435 105.235 30.825 105.525 ;
        RECT 35.705 105.375 102.905 105.625 ;
        RECT 35.705 105.355 71.615 105.375 ;
        RECT 107.125 105.255 113.515 105.545 ;
        RECT 23.850 104.655 34.355 104.990 ;
        RECT 59.325 104.790 69.875 105.125 ;
        RECT 106.540 104.675 117.020 105.010 ;
        RECT 23.200 104.070 26.120 104.370 ;
        RECT 29.665 104.055 33.035 104.355 ;
        RECT 37.915 104.150 39.220 104.530 ;
        RECT 39.920 104.150 43.220 104.530 ;
        RECT 43.920 104.150 47.220 104.530 ;
        RECT 47.920 104.150 49.280 104.530 ;
        RECT 51.255 104.150 52.720 104.530 ;
        RECT 53.420 104.150 56.720 104.530 ;
        RECT 57.420 104.150 60.720 104.530 ;
        RECT 61.420 104.150 62.600 104.530 ;
        RECT 76.510 104.170 77.815 104.550 ;
        RECT 82.515 104.170 85.815 104.550 ;
        RECT 86.515 104.170 87.875 104.550 ;
        RECT 89.850 104.170 91.315 104.550 ;
        RECT 92.015 104.170 95.315 104.550 ;
        RECT 100.015 104.170 101.195 104.550 ;
        RECT 39.380 103.805 39.760 103.840 ;
        RECT 21.415 103.320 21.795 103.700 ;
        RECT 23.820 103.335 25.600 103.625 ;
        RECT 27.075 103.425 28.265 103.710 ;
        RECT 31.195 103.305 32.505 103.625 ;
        RECT 39.115 103.495 42.125 103.805 ;
        RECT 39.380 103.460 39.760 103.495 ;
        RECT 43.380 103.460 44.470 103.840 ;
        RECT 47.380 103.835 47.760 103.840 ;
        RECT 44.900 103.470 47.765 103.835 ;
        RECT 52.880 103.815 53.260 103.840 ;
        RECT 52.865 103.495 55.010 103.815 ;
        RECT 47.380 103.460 47.760 103.470 ;
        RECT 52.880 103.460 53.260 103.495 ;
        RECT 55.925 103.460 57.260 103.840 ;
        RECT 60.880 103.820 61.260 103.840 ;
        RECT 77.975 103.825 78.355 103.860 ;
        RECT 58.415 103.500 61.325 103.820 ;
        RECT 77.710 103.515 80.720 103.825 ;
        RECT 60.880 103.460 61.260 103.500 ;
        RECT 77.975 103.480 78.355 103.515 ;
        RECT 81.975 103.480 83.065 103.860 ;
        RECT 85.975 103.855 86.355 103.860 ;
        RECT 83.495 103.490 86.360 103.855 ;
        RECT 91.475 103.835 91.855 103.860 ;
        RECT 91.460 103.515 93.605 103.835 ;
        RECT 85.975 103.480 86.355 103.490 ;
        RECT 91.475 103.480 91.855 103.515 ;
        RECT 94.520 103.480 95.855 103.860 ;
        RECT 99.475 103.840 99.855 103.860 ;
        RECT 97.010 103.520 99.920 103.840 ;
        RECT 99.475 103.480 99.855 103.520 ;
        RECT 104.105 103.340 104.485 103.720 ;
        RECT 106.510 103.355 108.290 103.645 ;
        RECT 109.765 103.445 110.955 103.730 ;
        RECT 113.885 103.325 115.195 103.645 ;
        RECT 22.550 102.720 22.930 103.100 ;
        RECT 26.295 102.760 26.675 103.140 ;
        RECT 29.005 102.750 29.385 103.130 ;
        RECT 30.415 102.595 33.595 102.915 ;
        RECT 105.240 102.740 105.620 103.120 ;
        RECT 108.985 102.780 109.365 103.160 ;
        RECT 111.695 102.770 112.075 103.150 ;
        RECT 113.105 102.615 116.285 102.935 ;
        RECT 37.730 102.150 39.220 102.530 ;
        RECT 39.920 102.150 41.205 102.530 ;
        RECT 59.235 102.150 60.720 102.530 ;
        RECT 61.420 102.150 62.495 102.530 ;
        RECT 76.325 102.170 77.815 102.550 ;
        RECT 100.015 102.170 101.090 102.550 ;
        RECT 39.380 101.460 40.470 101.840 ;
        RECT 41.425 101.470 42.945 101.830 ;
        RECT 43.865 101.465 56.715 101.800 ;
        RECT 60.880 101.795 61.260 101.840 ;
        RECT 60.145 101.495 61.455 101.795 ;
        RECT 60.880 101.460 61.260 101.495 ;
        RECT 77.975 101.480 79.065 101.860 ;
        RECT 80.020 101.490 81.540 101.850 ;
        RECT 82.460 101.485 95.310 101.820 ;
        RECT 99.475 101.815 99.855 101.860 ;
        RECT 98.740 101.515 100.050 101.815 ;
        RECT 99.475 101.480 99.855 101.515 ;
        RECT 68.535 100.950 101.485 100.985 ;
        RECT 36.235 100.620 101.485 100.950 ;
        RECT 36.235 100.600 69.315 100.620 ;
        RECT 103.280 100.610 107.540 100.965 ;
        RECT 101.485 100.025 107.130 100.030 ;
        RECT 117.745 100.025 118.125 105.855 ;
        RECT 126.625 105.805 131.125 106.115 ;
        RECT 202.875 105.835 207.005 106.135 ;
        RECT 122.585 105.255 128.975 105.545 ;
        RECT 122.000 104.675 138.020 105.010 ;
        RECT 186.800 104.775 192.715 105.110 ;
        RECT 190.070 104.755 192.715 104.775 ;
        RECT 121.350 104.090 124.270 104.390 ;
        RECT 127.815 104.075 131.185 104.375 ;
        RECT 167.395 104.135 170.695 104.515 ;
        RECT 171.395 104.135 174.695 104.515 ;
        RECT 180.895 104.135 184.195 104.515 ;
        RECT 184.895 104.135 188.195 104.515 ;
        RECT 119.565 103.340 119.945 103.720 ;
        RECT 121.970 103.355 123.750 103.645 ;
        RECT 125.225 103.445 126.415 103.730 ;
        RECT 129.345 103.325 130.655 103.645 ;
        RECT 120.700 102.740 121.080 103.120 ;
        RECT 124.445 102.780 124.825 103.160 ;
        RECT 127.155 102.770 127.535 103.150 ;
        RECT 128.565 102.615 131.745 102.935 ;
        RECT 167.395 102.135 168.680 102.515 ;
        RECT 186.710 102.135 188.195 102.515 ;
        RECT 118.845 101.530 122.995 101.800 ;
        RECT 168.900 101.455 170.420 101.815 ;
        RECT 118.495 100.025 122.590 100.030 ;
        RECT 74.830 100.020 107.130 100.025 ;
        RECT 117.375 100.020 122.590 100.025 ;
        RECT 20.345 100.005 24.440 100.010 ;
        RECT 74.830 100.005 132.405 100.020 ;
        RECT 200.500 100.005 200.880 105.835 ;
        RECT 209.380 105.785 213.880 106.095 ;
        RECT 218.335 105.835 222.465 106.135 ;
        RECT 205.340 105.235 211.730 105.525 ;
        RECT 204.755 104.655 215.410 104.990 ;
        RECT 204.105 104.070 207.025 104.370 ;
        RECT 210.570 104.055 213.940 104.355 ;
        RECT 202.320 103.320 202.700 103.700 ;
        RECT 204.725 103.335 206.505 103.625 ;
        RECT 207.980 103.425 209.170 103.710 ;
        RECT 212.100 103.305 213.410 103.625 ;
        RECT 203.455 102.720 203.835 103.100 ;
        RECT 207.200 102.760 207.580 103.140 ;
        RECT 209.910 102.750 210.290 103.130 ;
        RECT 211.320 102.595 214.500 102.915 ;
        RECT 201.250 100.005 205.345 100.010 ;
        RECT 215.960 100.005 216.340 105.835 ;
        RECT 224.840 105.785 229.340 106.095 ;
        RECT 316.485 105.855 320.615 106.155 ;
        RECT 267.525 105.625 299.270 105.645 ;
        RECT 220.800 105.235 227.190 105.525 ;
        RECT 232.070 105.375 299.270 105.625 ;
        RECT 232.070 105.355 267.980 105.375 ;
        RECT 303.490 105.255 309.880 105.545 ;
        RECT 220.215 104.655 230.720 104.990 ;
        RECT 255.690 104.790 266.240 105.125 ;
        RECT 302.905 104.675 313.385 105.010 ;
        RECT 219.565 104.070 222.485 104.370 ;
        RECT 226.030 104.055 229.400 104.355 ;
        RECT 234.280 104.150 235.585 104.530 ;
        RECT 236.285 104.150 239.585 104.530 ;
        RECT 240.285 104.150 243.585 104.530 ;
        RECT 244.285 104.150 245.645 104.530 ;
        RECT 247.620 104.150 249.085 104.530 ;
        RECT 249.785 104.150 253.085 104.530 ;
        RECT 253.785 104.150 257.085 104.530 ;
        RECT 257.785 104.150 258.965 104.530 ;
        RECT 272.875 104.170 274.180 104.550 ;
        RECT 278.880 104.170 282.180 104.550 ;
        RECT 282.880 104.170 284.240 104.550 ;
        RECT 286.215 104.170 287.680 104.550 ;
        RECT 288.380 104.170 291.680 104.550 ;
        RECT 296.380 104.170 297.560 104.550 ;
        RECT 235.745 103.805 236.125 103.840 ;
        RECT 217.780 103.320 218.160 103.700 ;
        RECT 220.185 103.335 221.965 103.625 ;
        RECT 223.440 103.425 224.630 103.710 ;
        RECT 227.560 103.305 228.870 103.625 ;
        RECT 235.480 103.495 238.490 103.805 ;
        RECT 235.745 103.460 236.125 103.495 ;
        RECT 239.745 103.460 240.835 103.840 ;
        RECT 243.745 103.835 244.125 103.840 ;
        RECT 241.265 103.470 244.130 103.835 ;
        RECT 249.245 103.815 249.625 103.840 ;
        RECT 249.230 103.495 251.375 103.815 ;
        RECT 243.745 103.460 244.125 103.470 ;
        RECT 249.245 103.460 249.625 103.495 ;
        RECT 252.290 103.460 253.625 103.840 ;
        RECT 257.245 103.820 257.625 103.840 ;
        RECT 274.340 103.825 274.720 103.860 ;
        RECT 254.780 103.500 257.690 103.820 ;
        RECT 274.075 103.515 277.085 103.825 ;
        RECT 257.245 103.460 257.625 103.500 ;
        RECT 274.340 103.480 274.720 103.515 ;
        RECT 278.340 103.480 279.430 103.860 ;
        RECT 282.340 103.855 282.720 103.860 ;
        RECT 279.860 103.490 282.725 103.855 ;
        RECT 287.840 103.835 288.220 103.860 ;
        RECT 287.825 103.515 289.970 103.835 ;
        RECT 282.340 103.480 282.720 103.490 ;
        RECT 287.840 103.480 288.220 103.515 ;
        RECT 290.885 103.480 292.220 103.860 ;
        RECT 295.840 103.840 296.220 103.860 ;
        RECT 293.375 103.520 296.285 103.840 ;
        RECT 295.840 103.480 296.220 103.520 ;
        RECT 300.470 103.340 300.850 103.720 ;
        RECT 302.875 103.355 304.655 103.645 ;
        RECT 306.130 103.445 307.320 103.730 ;
        RECT 310.250 103.325 311.560 103.645 ;
        RECT 218.915 102.720 219.295 103.100 ;
        RECT 222.660 102.760 223.040 103.140 ;
        RECT 225.370 102.750 225.750 103.130 ;
        RECT 226.780 102.595 229.960 102.915 ;
        RECT 301.605 102.740 301.985 103.120 ;
        RECT 305.350 102.780 305.730 103.160 ;
        RECT 308.060 102.770 308.440 103.150 ;
        RECT 309.470 102.615 312.650 102.935 ;
        RECT 234.095 102.150 235.585 102.530 ;
        RECT 236.285 102.150 237.570 102.530 ;
        RECT 255.600 102.150 257.085 102.530 ;
        RECT 257.785 102.150 258.860 102.530 ;
        RECT 272.690 102.170 274.180 102.550 ;
        RECT 296.380 102.170 297.455 102.550 ;
        RECT 235.745 101.460 236.835 101.840 ;
        RECT 237.790 101.470 239.310 101.830 ;
        RECT 240.230 101.465 253.080 101.800 ;
        RECT 257.245 101.795 257.625 101.840 ;
        RECT 256.510 101.495 257.820 101.795 ;
        RECT 257.245 101.460 257.625 101.495 ;
        RECT 274.340 101.480 275.430 101.860 ;
        RECT 276.385 101.490 277.905 101.850 ;
        RECT 278.825 101.485 291.675 101.820 ;
        RECT 295.840 101.815 296.220 101.860 ;
        RECT 295.105 101.515 296.415 101.815 ;
        RECT 295.840 101.480 296.220 101.515 ;
        RECT 264.900 100.950 297.850 100.985 ;
        RECT 232.600 100.620 297.850 100.950 ;
        RECT 232.600 100.600 265.680 100.620 ;
        RECT 299.645 100.610 303.905 100.965 ;
        RECT 297.850 100.025 303.495 100.030 ;
        RECT 314.110 100.025 314.490 105.855 ;
        RECT 322.990 105.805 327.490 106.115 ;
        RECT 399.275 105.785 403.405 106.085 ;
        RECT 318.950 105.255 325.340 105.545 ;
        RECT 318.365 104.675 334.385 105.010 ;
        RECT 383.190 104.735 389.105 105.070 ;
        RECT 386.460 104.715 389.105 104.735 ;
        RECT 317.715 104.090 320.635 104.390 ;
        RECT 324.180 104.075 327.550 104.375 ;
        RECT 363.785 104.095 367.085 104.475 ;
        RECT 367.785 104.095 371.085 104.475 ;
        RECT 377.285 104.095 380.585 104.475 ;
        RECT 381.285 104.095 384.585 104.475 ;
        RECT 315.930 103.340 316.310 103.720 ;
        RECT 318.335 103.355 320.115 103.645 ;
        RECT 321.590 103.445 322.780 103.730 ;
        RECT 325.710 103.325 327.020 103.645 ;
        RECT 317.065 102.740 317.445 103.120 ;
        RECT 320.810 102.780 321.190 103.160 ;
        RECT 323.520 102.770 323.900 103.150 ;
        RECT 324.930 102.615 328.110 102.935 ;
        RECT 363.785 102.095 365.070 102.475 ;
        RECT 383.100 102.095 384.585 102.475 ;
        RECT 315.210 101.530 319.360 101.800 ;
        RECT 365.290 101.415 366.810 101.775 ;
        RECT 314.860 100.025 318.955 100.030 ;
        RECT 271.195 100.020 303.495 100.025 ;
        RECT 313.740 100.020 318.955 100.025 ;
        RECT 216.710 100.005 220.805 100.010 ;
        RECT 271.195 100.005 328.770 100.020 ;
        RECT 3.765 100.000 8.980 100.005 ;
        RECT 19.225 100.000 24.440 100.005 ;
        RECT 34.685 100.000 132.405 100.005 ;
        RECT -82.785 99.000 -56.130 99.900 ;
        RECT -32.460 99.080 -5.805 99.980 ;
        RECT 3.765 99.125 132.405 100.000 ;
        RECT 200.130 100.000 205.345 100.005 ;
        RECT 215.590 100.000 220.805 100.005 ;
        RECT 231.050 100.000 328.770 100.005 ;
        RECT 3.765 99.105 74.935 99.125 ;
        RECT 163.710 99.090 190.365 99.990 ;
        RECT 200.130 99.125 328.770 100.000 ;
        RECT 396.900 99.955 397.280 105.785 ;
        RECT 405.780 105.735 410.280 106.045 ;
        RECT 414.735 105.785 418.865 106.085 ;
        RECT 401.740 105.185 408.130 105.475 ;
        RECT 401.155 104.605 411.810 104.940 ;
        RECT 400.505 104.020 403.425 104.320 ;
        RECT 406.970 104.005 410.340 104.305 ;
        RECT 398.720 103.270 399.100 103.650 ;
        RECT 401.125 103.285 402.905 103.575 ;
        RECT 404.380 103.375 405.570 103.660 ;
        RECT 408.500 103.255 409.810 103.575 ;
        RECT 399.855 102.670 400.235 103.050 ;
        RECT 403.600 102.710 403.980 103.090 ;
        RECT 406.310 102.700 406.690 103.080 ;
        RECT 407.720 102.545 410.900 102.865 ;
        RECT 397.650 99.955 401.745 99.960 ;
        RECT 412.360 99.955 412.740 105.785 ;
        RECT 421.240 105.735 425.740 106.045 ;
        RECT 512.885 105.805 517.015 106.105 ;
        RECT 463.925 105.575 495.670 105.595 ;
        RECT 417.200 105.185 423.590 105.475 ;
        RECT 428.470 105.325 495.670 105.575 ;
        RECT 428.470 105.305 464.380 105.325 ;
        RECT 499.890 105.205 506.280 105.495 ;
        RECT 416.615 104.605 427.120 104.940 ;
        RECT 452.090 104.740 462.640 105.075 ;
        RECT 499.305 104.625 509.785 104.960 ;
        RECT 415.965 104.020 418.885 104.320 ;
        RECT 422.430 104.005 425.800 104.305 ;
        RECT 430.680 104.100 431.985 104.480 ;
        RECT 432.685 104.100 435.985 104.480 ;
        RECT 436.685 104.100 439.985 104.480 ;
        RECT 440.685 104.100 442.045 104.480 ;
        RECT 444.020 104.100 445.485 104.480 ;
        RECT 446.185 104.100 449.485 104.480 ;
        RECT 450.185 104.100 453.485 104.480 ;
        RECT 454.185 104.100 455.365 104.480 ;
        RECT 469.275 104.120 470.580 104.500 ;
        RECT 475.280 104.120 478.580 104.500 ;
        RECT 479.280 104.120 480.640 104.500 ;
        RECT 482.615 104.120 484.080 104.500 ;
        RECT 484.780 104.120 488.080 104.500 ;
        RECT 492.780 104.120 493.960 104.500 ;
        RECT 432.145 103.755 432.525 103.790 ;
        RECT 414.180 103.270 414.560 103.650 ;
        RECT 416.585 103.285 418.365 103.575 ;
        RECT 419.840 103.375 421.030 103.660 ;
        RECT 423.960 103.255 425.270 103.575 ;
        RECT 431.880 103.445 434.890 103.755 ;
        RECT 432.145 103.410 432.525 103.445 ;
        RECT 436.145 103.410 437.235 103.790 ;
        RECT 440.145 103.785 440.525 103.790 ;
        RECT 437.665 103.420 440.530 103.785 ;
        RECT 445.645 103.765 446.025 103.790 ;
        RECT 445.630 103.445 447.775 103.765 ;
        RECT 440.145 103.410 440.525 103.420 ;
        RECT 445.645 103.410 446.025 103.445 ;
        RECT 448.690 103.410 450.025 103.790 ;
        RECT 453.645 103.770 454.025 103.790 ;
        RECT 470.740 103.775 471.120 103.810 ;
        RECT 451.180 103.450 454.090 103.770 ;
        RECT 470.475 103.465 473.485 103.775 ;
        RECT 453.645 103.410 454.025 103.450 ;
        RECT 470.740 103.430 471.120 103.465 ;
        RECT 474.740 103.430 475.830 103.810 ;
        RECT 478.740 103.805 479.120 103.810 ;
        RECT 476.260 103.440 479.125 103.805 ;
        RECT 484.240 103.785 484.620 103.810 ;
        RECT 484.225 103.465 486.370 103.785 ;
        RECT 478.740 103.430 479.120 103.440 ;
        RECT 484.240 103.430 484.620 103.465 ;
        RECT 487.285 103.430 488.620 103.810 ;
        RECT 492.240 103.790 492.620 103.810 ;
        RECT 489.775 103.470 492.685 103.790 ;
        RECT 492.240 103.430 492.620 103.470 ;
        RECT 496.870 103.290 497.250 103.670 ;
        RECT 499.275 103.305 501.055 103.595 ;
        RECT 502.530 103.395 503.720 103.680 ;
        RECT 506.650 103.275 507.960 103.595 ;
        RECT 415.315 102.670 415.695 103.050 ;
        RECT 419.060 102.710 419.440 103.090 ;
        RECT 421.770 102.700 422.150 103.080 ;
        RECT 423.180 102.545 426.360 102.865 ;
        RECT 498.005 102.690 498.385 103.070 ;
        RECT 501.750 102.730 502.130 103.110 ;
        RECT 504.460 102.720 504.840 103.100 ;
        RECT 505.870 102.565 509.050 102.885 ;
        RECT 430.495 102.100 431.985 102.480 ;
        RECT 432.685 102.100 433.970 102.480 ;
        RECT 452.000 102.100 453.485 102.480 ;
        RECT 454.185 102.100 455.260 102.480 ;
        RECT 469.090 102.120 470.580 102.500 ;
        RECT 492.780 102.120 493.855 102.500 ;
        RECT 432.145 101.410 433.235 101.790 ;
        RECT 434.190 101.420 435.710 101.780 ;
        RECT 436.630 101.415 449.480 101.750 ;
        RECT 453.645 101.745 454.025 101.790 ;
        RECT 452.910 101.445 454.220 101.745 ;
        RECT 453.645 101.410 454.025 101.445 ;
        RECT 470.740 101.430 471.830 101.810 ;
        RECT 472.785 101.440 474.305 101.800 ;
        RECT 475.225 101.435 488.075 101.770 ;
        RECT 492.240 101.765 492.620 101.810 ;
        RECT 491.505 101.465 492.815 101.765 ;
        RECT 492.240 101.430 492.620 101.465 ;
        RECT 461.300 100.900 494.250 100.935 ;
        RECT 429.000 100.570 494.250 100.900 ;
        RECT 429.000 100.550 462.080 100.570 ;
        RECT 496.045 100.560 500.305 100.915 ;
        RECT 494.250 99.975 499.895 99.980 ;
        RECT 510.510 99.975 510.890 105.805 ;
        RECT 519.390 105.755 523.890 106.065 ;
        RECT 595.650 105.820 599.780 106.120 ;
        RECT 515.350 105.205 521.740 105.495 ;
        RECT 514.765 104.625 530.785 104.960 ;
        RECT 579.510 104.780 585.425 105.115 ;
        RECT 582.780 104.760 585.425 104.780 ;
        RECT 514.115 104.040 517.035 104.340 ;
        RECT 520.580 104.025 523.950 104.325 ;
        RECT 560.105 104.140 563.405 104.520 ;
        RECT 564.105 104.140 567.405 104.520 ;
        RECT 573.605 104.140 576.905 104.520 ;
        RECT 577.605 104.140 580.905 104.520 ;
        RECT 512.330 103.290 512.710 103.670 ;
        RECT 514.735 103.305 516.515 103.595 ;
        RECT 517.990 103.395 519.180 103.680 ;
        RECT 522.110 103.275 523.420 103.595 ;
        RECT 513.465 102.690 513.845 103.070 ;
        RECT 517.210 102.730 517.590 103.110 ;
        RECT 519.920 102.720 520.300 103.100 ;
        RECT 521.330 102.565 524.510 102.885 ;
        RECT 560.105 102.140 561.390 102.520 ;
        RECT 579.420 102.140 580.905 102.520 ;
        RECT 511.610 101.480 515.760 101.750 ;
        RECT 561.610 101.460 563.130 101.820 ;
        RECT 511.260 99.975 515.355 99.980 ;
        RECT 467.595 99.970 499.895 99.975 ;
        RECT 510.140 99.970 515.355 99.975 ;
        RECT 413.110 99.955 417.205 99.960 ;
        RECT 467.595 99.955 525.170 99.970 ;
        RECT 396.530 99.950 401.745 99.955 ;
        RECT 411.990 99.950 417.205 99.955 ;
        RECT 427.450 99.950 525.170 99.955 ;
        RECT 200.130 99.105 271.300 99.125 ;
        RECT 360.100 99.050 386.755 99.950 ;
        RECT 396.530 99.075 525.170 99.950 ;
        RECT 556.420 99.095 583.075 99.995 ;
        RECT 593.275 99.990 593.655 105.820 ;
        RECT 602.155 105.770 606.655 106.080 ;
        RECT 611.110 105.820 615.240 106.120 ;
        RECT 598.115 105.220 604.505 105.510 ;
        RECT 597.530 104.640 608.185 104.975 ;
        RECT 596.880 104.055 599.800 104.355 ;
        RECT 603.345 104.040 606.715 104.340 ;
        RECT 595.095 103.305 595.475 103.685 ;
        RECT 597.500 103.320 599.280 103.610 ;
        RECT 600.755 103.410 601.945 103.695 ;
        RECT 604.875 103.290 606.185 103.610 ;
        RECT 596.230 102.705 596.610 103.085 ;
        RECT 599.975 102.745 600.355 103.125 ;
        RECT 602.685 102.735 603.065 103.115 ;
        RECT 604.095 102.580 607.275 102.900 ;
        RECT 594.025 99.990 598.120 99.995 ;
        RECT 608.735 99.990 609.115 105.820 ;
        RECT 617.615 105.770 622.115 106.080 ;
        RECT 709.260 105.840 713.390 106.140 ;
        RECT 660.300 105.610 692.045 105.630 ;
        RECT 613.575 105.220 619.965 105.510 ;
        RECT 624.845 105.360 692.045 105.610 ;
        RECT 624.845 105.340 660.755 105.360 ;
        RECT 696.265 105.240 702.655 105.530 ;
        RECT 612.990 104.640 623.495 104.975 ;
        RECT 648.465 104.775 659.015 105.110 ;
        RECT 695.680 104.660 706.160 104.995 ;
        RECT 612.340 104.055 615.260 104.355 ;
        RECT 618.805 104.040 622.175 104.340 ;
        RECT 627.055 104.135 628.360 104.515 ;
        RECT 629.060 104.135 632.360 104.515 ;
        RECT 633.060 104.135 636.360 104.515 ;
        RECT 637.060 104.135 638.420 104.515 ;
        RECT 640.395 104.135 641.860 104.515 ;
        RECT 642.560 104.135 645.860 104.515 ;
        RECT 646.560 104.135 649.860 104.515 ;
        RECT 650.560 104.135 651.740 104.515 ;
        RECT 665.650 104.155 666.955 104.535 ;
        RECT 671.655 104.155 674.955 104.535 ;
        RECT 675.655 104.155 677.015 104.535 ;
        RECT 678.990 104.155 680.455 104.535 ;
        RECT 681.155 104.155 684.455 104.535 ;
        RECT 689.155 104.155 690.335 104.535 ;
        RECT 628.520 103.790 628.900 103.825 ;
        RECT 610.555 103.305 610.935 103.685 ;
        RECT 612.960 103.320 614.740 103.610 ;
        RECT 616.215 103.410 617.405 103.695 ;
        RECT 620.335 103.290 621.645 103.610 ;
        RECT 628.255 103.480 631.265 103.790 ;
        RECT 628.520 103.445 628.900 103.480 ;
        RECT 632.520 103.445 633.610 103.825 ;
        RECT 636.520 103.820 636.900 103.825 ;
        RECT 634.040 103.455 636.905 103.820 ;
        RECT 642.020 103.800 642.400 103.825 ;
        RECT 642.005 103.480 644.150 103.800 ;
        RECT 636.520 103.445 636.900 103.455 ;
        RECT 642.020 103.445 642.400 103.480 ;
        RECT 645.065 103.445 646.400 103.825 ;
        RECT 650.020 103.805 650.400 103.825 ;
        RECT 667.115 103.810 667.495 103.845 ;
        RECT 647.555 103.485 650.465 103.805 ;
        RECT 666.850 103.500 669.860 103.810 ;
        RECT 650.020 103.445 650.400 103.485 ;
        RECT 667.115 103.465 667.495 103.500 ;
        RECT 671.115 103.465 672.205 103.845 ;
        RECT 675.115 103.840 675.495 103.845 ;
        RECT 672.635 103.475 675.500 103.840 ;
        RECT 680.615 103.820 680.995 103.845 ;
        RECT 680.600 103.500 682.745 103.820 ;
        RECT 675.115 103.465 675.495 103.475 ;
        RECT 680.615 103.465 680.995 103.500 ;
        RECT 683.660 103.465 684.995 103.845 ;
        RECT 688.615 103.825 688.995 103.845 ;
        RECT 686.150 103.505 689.060 103.825 ;
        RECT 688.615 103.465 688.995 103.505 ;
        RECT 693.245 103.325 693.625 103.705 ;
        RECT 695.650 103.340 697.430 103.630 ;
        RECT 698.905 103.430 700.095 103.715 ;
        RECT 703.025 103.310 704.335 103.630 ;
        RECT 611.690 102.705 612.070 103.085 ;
        RECT 615.435 102.745 615.815 103.125 ;
        RECT 618.145 102.735 618.525 103.115 ;
        RECT 619.555 102.580 622.735 102.900 ;
        RECT 694.380 102.725 694.760 103.105 ;
        RECT 698.125 102.765 698.505 103.145 ;
        RECT 700.835 102.755 701.215 103.135 ;
        RECT 702.245 102.600 705.425 102.920 ;
        RECT 626.870 102.135 628.360 102.515 ;
        RECT 629.060 102.135 630.345 102.515 ;
        RECT 648.375 102.135 649.860 102.515 ;
        RECT 650.560 102.135 651.635 102.515 ;
        RECT 665.465 102.155 666.955 102.535 ;
        RECT 689.155 102.155 690.230 102.535 ;
        RECT 628.520 101.445 629.610 101.825 ;
        RECT 630.565 101.455 632.085 101.815 ;
        RECT 633.005 101.450 645.855 101.785 ;
        RECT 650.020 101.780 650.400 101.825 ;
        RECT 649.285 101.480 650.595 101.780 ;
        RECT 650.020 101.445 650.400 101.480 ;
        RECT 667.115 101.465 668.205 101.845 ;
        RECT 669.160 101.475 670.680 101.835 ;
        RECT 671.600 101.470 684.450 101.805 ;
        RECT 688.615 101.800 688.995 101.845 ;
        RECT 687.880 101.500 689.190 101.800 ;
        RECT 688.615 101.465 688.995 101.500 ;
        RECT 657.675 100.935 690.625 100.970 ;
        RECT 625.375 100.605 690.625 100.935 ;
        RECT 625.375 100.585 658.455 100.605 ;
        RECT 692.420 100.595 696.680 100.950 ;
        RECT 690.625 100.010 696.270 100.015 ;
        RECT 706.885 100.010 707.265 105.840 ;
        RECT 715.765 105.790 720.265 106.100 ;
        RECT 791.990 105.820 796.120 106.120 ;
        RECT 711.725 105.240 718.115 105.530 ;
        RECT 711.140 104.660 727.160 104.995 ;
        RECT 775.875 104.785 781.790 105.120 ;
        RECT 779.145 104.765 781.790 104.785 ;
        RECT 710.490 104.075 713.410 104.375 ;
        RECT 716.955 104.060 720.325 104.360 ;
        RECT 756.470 104.145 759.770 104.525 ;
        RECT 760.470 104.145 763.770 104.525 ;
        RECT 769.970 104.145 773.270 104.525 ;
        RECT 773.970 104.145 777.270 104.525 ;
        RECT 708.705 103.325 709.085 103.705 ;
        RECT 711.110 103.340 712.890 103.630 ;
        RECT 714.365 103.430 715.555 103.715 ;
        RECT 718.485 103.310 719.795 103.630 ;
        RECT 709.840 102.725 710.220 103.105 ;
        RECT 713.585 102.765 713.965 103.145 ;
        RECT 716.295 102.755 716.675 103.135 ;
        RECT 717.705 102.600 720.885 102.920 ;
        RECT 756.470 102.145 757.755 102.525 ;
        RECT 775.785 102.145 777.270 102.525 ;
        RECT 707.985 101.515 712.135 101.785 ;
        RECT 757.975 101.465 759.495 101.825 ;
        RECT 707.635 100.010 711.730 100.015 ;
        RECT 663.970 100.005 696.270 100.010 ;
        RECT 706.515 100.005 711.730 100.010 ;
        RECT 609.485 99.990 613.580 99.995 ;
        RECT 663.970 99.990 721.545 100.005 ;
        RECT 592.905 99.985 598.120 99.990 ;
        RECT 608.365 99.985 613.580 99.990 ;
        RECT 623.825 99.985 721.545 99.990 ;
        RECT 592.905 99.110 721.545 99.985 ;
        RECT 592.905 99.090 664.075 99.110 ;
        RECT 752.785 99.100 779.440 100.000 ;
        RECT 789.615 99.990 789.995 105.820 ;
        RECT 798.495 105.770 802.995 106.080 ;
        RECT 807.450 105.820 811.580 106.120 ;
        RECT 794.455 105.220 800.845 105.510 ;
        RECT 793.870 104.640 804.525 104.975 ;
        RECT 793.220 104.055 796.140 104.355 ;
        RECT 799.685 104.040 803.055 104.340 ;
        RECT 791.435 103.305 791.815 103.685 ;
        RECT 793.840 103.320 795.620 103.610 ;
        RECT 797.095 103.410 798.285 103.695 ;
        RECT 801.215 103.290 802.525 103.610 ;
        RECT 792.570 102.705 792.950 103.085 ;
        RECT 796.315 102.745 796.695 103.125 ;
        RECT 799.025 102.735 799.405 103.115 ;
        RECT 800.435 102.580 803.615 102.900 ;
        RECT 790.365 99.990 794.460 99.995 ;
        RECT 805.075 99.990 805.455 105.820 ;
        RECT 813.955 105.770 818.455 106.080 ;
        RECT 905.600 105.840 909.730 106.140 ;
        RECT 856.640 105.610 888.385 105.630 ;
        RECT 809.915 105.220 816.305 105.510 ;
        RECT 821.185 105.360 888.385 105.610 ;
        RECT 821.185 105.340 857.095 105.360 ;
        RECT 892.605 105.240 898.995 105.530 ;
        RECT 809.330 104.640 819.835 104.975 ;
        RECT 844.805 104.775 855.355 105.110 ;
        RECT 892.020 104.660 902.500 104.995 ;
        RECT 808.680 104.055 811.600 104.355 ;
        RECT 815.145 104.040 818.515 104.340 ;
        RECT 823.395 104.135 824.700 104.515 ;
        RECT 825.400 104.135 828.700 104.515 ;
        RECT 829.400 104.135 832.700 104.515 ;
        RECT 833.400 104.135 834.760 104.515 ;
        RECT 836.735 104.135 838.200 104.515 ;
        RECT 838.900 104.135 842.200 104.515 ;
        RECT 842.900 104.135 846.200 104.515 ;
        RECT 846.900 104.135 848.080 104.515 ;
        RECT 861.990 104.155 863.295 104.535 ;
        RECT 867.995 104.155 871.295 104.535 ;
        RECT 871.995 104.155 873.355 104.535 ;
        RECT 875.330 104.155 876.795 104.535 ;
        RECT 877.495 104.155 880.795 104.535 ;
        RECT 885.495 104.155 886.675 104.535 ;
        RECT 824.860 103.790 825.240 103.825 ;
        RECT 806.895 103.305 807.275 103.685 ;
        RECT 809.300 103.320 811.080 103.610 ;
        RECT 812.555 103.410 813.745 103.695 ;
        RECT 816.675 103.290 817.985 103.610 ;
        RECT 824.595 103.480 827.605 103.790 ;
        RECT 824.860 103.445 825.240 103.480 ;
        RECT 828.860 103.445 829.950 103.825 ;
        RECT 832.860 103.820 833.240 103.825 ;
        RECT 830.380 103.455 833.245 103.820 ;
        RECT 838.360 103.800 838.740 103.825 ;
        RECT 838.345 103.480 840.490 103.800 ;
        RECT 832.860 103.445 833.240 103.455 ;
        RECT 838.360 103.445 838.740 103.480 ;
        RECT 841.405 103.445 842.740 103.825 ;
        RECT 846.360 103.805 846.740 103.825 ;
        RECT 863.455 103.810 863.835 103.845 ;
        RECT 843.895 103.485 846.805 103.805 ;
        RECT 863.190 103.500 866.200 103.810 ;
        RECT 846.360 103.445 846.740 103.485 ;
        RECT 863.455 103.465 863.835 103.500 ;
        RECT 867.455 103.465 868.545 103.845 ;
        RECT 871.455 103.840 871.835 103.845 ;
        RECT 868.975 103.475 871.840 103.840 ;
        RECT 876.955 103.820 877.335 103.845 ;
        RECT 876.940 103.500 879.085 103.820 ;
        RECT 871.455 103.465 871.835 103.475 ;
        RECT 876.955 103.465 877.335 103.500 ;
        RECT 880.000 103.465 881.335 103.845 ;
        RECT 884.955 103.825 885.335 103.845 ;
        RECT 882.490 103.505 885.400 103.825 ;
        RECT 884.955 103.465 885.335 103.505 ;
        RECT 889.585 103.325 889.965 103.705 ;
        RECT 891.990 103.340 893.770 103.630 ;
        RECT 895.245 103.430 896.435 103.715 ;
        RECT 899.365 103.310 900.675 103.630 ;
        RECT 808.030 102.705 808.410 103.085 ;
        RECT 811.775 102.745 812.155 103.125 ;
        RECT 814.485 102.735 814.865 103.115 ;
        RECT 815.895 102.580 819.075 102.900 ;
        RECT 890.720 102.725 891.100 103.105 ;
        RECT 894.465 102.765 894.845 103.145 ;
        RECT 897.175 102.755 897.555 103.135 ;
        RECT 898.585 102.600 901.765 102.920 ;
        RECT 823.210 102.135 824.700 102.515 ;
        RECT 825.400 102.135 826.685 102.515 ;
        RECT 844.715 102.135 846.200 102.515 ;
        RECT 846.900 102.135 847.975 102.515 ;
        RECT 861.805 102.155 863.295 102.535 ;
        RECT 885.495 102.155 886.570 102.535 ;
        RECT 824.860 101.445 825.950 101.825 ;
        RECT 826.905 101.455 828.425 101.815 ;
        RECT 829.345 101.450 842.195 101.785 ;
        RECT 846.360 101.780 846.740 101.825 ;
        RECT 845.625 101.480 846.935 101.780 ;
        RECT 846.360 101.445 846.740 101.480 ;
        RECT 863.455 101.465 864.545 101.845 ;
        RECT 865.500 101.475 867.020 101.835 ;
        RECT 867.940 101.470 880.790 101.805 ;
        RECT 884.955 101.800 885.335 101.845 ;
        RECT 884.220 101.500 885.530 101.800 ;
        RECT 884.955 101.465 885.335 101.500 ;
        RECT 854.015 100.935 886.965 100.970 ;
        RECT 821.715 100.605 886.965 100.935 ;
        RECT 821.715 100.585 854.795 100.605 ;
        RECT 888.760 100.595 893.020 100.950 ;
        RECT 886.965 100.010 892.610 100.015 ;
        RECT 903.225 100.010 903.605 105.840 ;
        RECT 912.105 105.790 916.605 106.100 ;
        RECT 988.330 105.820 992.460 106.120 ;
        RECT 908.065 105.240 914.455 105.530 ;
        RECT 907.480 104.660 923.500 104.995 ;
        RECT 972.260 104.770 978.175 105.105 ;
        RECT 975.530 104.750 978.175 104.770 ;
        RECT 906.830 104.075 909.750 104.375 ;
        RECT 913.295 104.060 916.665 104.360 ;
        RECT 952.855 104.130 956.155 104.510 ;
        RECT 956.855 104.130 960.155 104.510 ;
        RECT 966.355 104.130 969.655 104.510 ;
        RECT 970.355 104.130 973.655 104.510 ;
        RECT 905.045 103.325 905.425 103.705 ;
        RECT 907.450 103.340 909.230 103.630 ;
        RECT 910.705 103.430 911.895 103.715 ;
        RECT 914.825 103.310 916.135 103.630 ;
        RECT 906.180 102.725 906.560 103.105 ;
        RECT 909.925 102.765 910.305 103.145 ;
        RECT 912.635 102.755 913.015 103.135 ;
        RECT 914.045 102.600 917.225 102.920 ;
        RECT 952.855 102.130 954.140 102.510 ;
        RECT 972.170 102.130 973.655 102.510 ;
        RECT 904.325 101.515 908.475 101.785 ;
        RECT 954.360 101.450 955.880 101.810 ;
        RECT 903.975 100.010 908.070 100.015 ;
        RECT 860.310 100.005 892.610 100.010 ;
        RECT 902.855 100.005 908.070 100.010 ;
        RECT 805.825 99.990 809.920 99.995 ;
        RECT 860.310 99.990 917.885 100.005 ;
        RECT 985.955 99.990 986.335 105.820 ;
        RECT 994.835 105.770 999.335 106.080 ;
        RECT 1003.790 105.820 1007.920 106.120 ;
        RECT 990.795 105.220 997.185 105.510 ;
        RECT 990.210 104.640 1000.865 104.975 ;
        RECT 989.560 104.055 992.480 104.355 ;
        RECT 996.025 104.040 999.395 104.340 ;
        RECT 987.775 103.305 988.155 103.685 ;
        RECT 990.180 103.320 991.960 103.610 ;
        RECT 993.435 103.410 994.625 103.695 ;
        RECT 997.555 103.290 998.865 103.610 ;
        RECT 988.910 102.705 989.290 103.085 ;
        RECT 992.655 102.745 993.035 103.125 ;
        RECT 995.365 102.735 995.745 103.115 ;
        RECT 996.775 102.580 999.955 102.900 ;
        RECT 986.705 99.990 990.800 99.995 ;
        RECT 1001.415 99.990 1001.795 105.820 ;
        RECT 1010.295 105.770 1014.795 106.080 ;
        RECT 1101.940 105.840 1106.070 106.140 ;
        RECT 1052.980 105.610 1084.725 105.630 ;
        RECT 1006.255 105.220 1012.645 105.510 ;
        RECT 1017.525 105.360 1084.725 105.610 ;
        RECT 1017.525 105.340 1053.435 105.360 ;
        RECT 1088.945 105.240 1095.335 105.530 ;
        RECT 1005.670 104.640 1016.175 104.975 ;
        RECT 1041.145 104.775 1051.695 105.110 ;
        RECT 1088.360 104.660 1098.840 104.995 ;
        RECT 1005.020 104.055 1007.940 104.355 ;
        RECT 1011.485 104.040 1014.855 104.340 ;
        RECT 1019.735 104.135 1021.040 104.515 ;
        RECT 1021.740 104.135 1025.040 104.515 ;
        RECT 1025.740 104.135 1029.040 104.515 ;
        RECT 1029.740 104.135 1031.100 104.515 ;
        RECT 1033.075 104.135 1034.540 104.515 ;
        RECT 1035.240 104.135 1038.540 104.515 ;
        RECT 1039.240 104.135 1042.540 104.515 ;
        RECT 1043.240 104.135 1044.420 104.515 ;
        RECT 1058.330 104.155 1059.635 104.535 ;
        RECT 1064.335 104.155 1067.635 104.535 ;
        RECT 1068.335 104.155 1069.695 104.535 ;
        RECT 1071.670 104.155 1073.135 104.535 ;
        RECT 1073.835 104.155 1077.135 104.535 ;
        RECT 1081.835 104.155 1083.015 104.535 ;
        RECT 1021.200 103.790 1021.580 103.825 ;
        RECT 1003.235 103.305 1003.615 103.685 ;
        RECT 1005.640 103.320 1007.420 103.610 ;
        RECT 1008.895 103.410 1010.085 103.695 ;
        RECT 1013.015 103.290 1014.325 103.610 ;
        RECT 1020.935 103.480 1023.945 103.790 ;
        RECT 1021.200 103.445 1021.580 103.480 ;
        RECT 1025.200 103.445 1026.290 103.825 ;
        RECT 1029.200 103.820 1029.580 103.825 ;
        RECT 1026.720 103.455 1029.585 103.820 ;
        RECT 1034.700 103.800 1035.080 103.825 ;
        RECT 1034.685 103.480 1036.830 103.800 ;
        RECT 1029.200 103.445 1029.580 103.455 ;
        RECT 1034.700 103.445 1035.080 103.480 ;
        RECT 1037.745 103.445 1039.080 103.825 ;
        RECT 1042.700 103.805 1043.080 103.825 ;
        RECT 1059.795 103.810 1060.175 103.845 ;
        RECT 1040.235 103.485 1043.145 103.805 ;
        RECT 1059.530 103.500 1062.540 103.810 ;
        RECT 1042.700 103.445 1043.080 103.485 ;
        RECT 1059.795 103.465 1060.175 103.500 ;
        RECT 1063.795 103.465 1064.885 103.845 ;
        RECT 1067.795 103.840 1068.175 103.845 ;
        RECT 1065.315 103.475 1068.180 103.840 ;
        RECT 1073.295 103.820 1073.675 103.845 ;
        RECT 1073.280 103.500 1075.425 103.820 ;
        RECT 1067.795 103.465 1068.175 103.475 ;
        RECT 1073.295 103.465 1073.675 103.500 ;
        RECT 1076.340 103.465 1077.675 103.845 ;
        RECT 1081.295 103.825 1081.675 103.845 ;
        RECT 1078.830 103.505 1081.740 103.825 ;
        RECT 1081.295 103.465 1081.675 103.505 ;
        RECT 1085.925 103.325 1086.305 103.705 ;
        RECT 1088.330 103.340 1090.110 103.630 ;
        RECT 1091.585 103.430 1092.775 103.715 ;
        RECT 1095.705 103.310 1097.015 103.630 ;
        RECT 1004.370 102.705 1004.750 103.085 ;
        RECT 1008.115 102.745 1008.495 103.125 ;
        RECT 1010.825 102.735 1011.205 103.115 ;
        RECT 1012.235 102.580 1015.415 102.900 ;
        RECT 1087.060 102.725 1087.440 103.105 ;
        RECT 1090.805 102.765 1091.185 103.145 ;
        RECT 1093.515 102.755 1093.895 103.135 ;
        RECT 1094.925 102.600 1098.105 102.920 ;
        RECT 1019.550 102.135 1021.040 102.515 ;
        RECT 1021.740 102.135 1023.025 102.515 ;
        RECT 1041.055 102.135 1042.540 102.515 ;
        RECT 1043.240 102.135 1044.315 102.515 ;
        RECT 1058.145 102.155 1059.635 102.535 ;
        RECT 1081.835 102.155 1082.910 102.535 ;
        RECT 1021.200 101.445 1022.290 101.825 ;
        RECT 1023.245 101.455 1024.765 101.815 ;
        RECT 1025.685 101.450 1038.535 101.785 ;
        RECT 1042.700 101.780 1043.080 101.825 ;
        RECT 1041.965 101.480 1043.275 101.780 ;
        RECT 1042.700 101.445 1043.080 101.480 ;
        RECT 1059.795 101.465 1060.885 101.845 ;
        RECT 1061.840 101.475 1063.360 101.835 ;
        RECT 1064.280 101.470 1077.130 101.805 ;
        RECT 1081.295 101.800 1081.675 101.845 ;
        RECT 1080.560 101.500 1081.870 101.800 ;
        RECT 1081.295 101.465 1081.675 101.500 ;
        RECT 1050.355 100.935 1083.305 100.970 ;
        RECT 1018.055 100.605 1083.305 100.935 ;
        RECT 1018.055 100.585 1051.135 100.605 ;
        RECT 1085.100 100.595 1089.360 100.950 ;
        RECT 1083.305 100.010 1088.950 100.015 ;
        RECT 1099.565 100.010 1099.945 105.840 ;
        RECT 1108.445 105.790 1112.945 106.100 ;
        RECT 1184.670 105.820 1188.800 106.120 ;
        RECT 1104.405 105.240 1110.795 105.530 ;
        RECT 1103.820 104.660 1119.840 104.995 ;
        RECT 1168.585 104.775 1174.500 105.110 ;
        RECT 1171.855 104.755 1174.500 104.775 ;
        RECT 1103.170 104.075 1106.090 104.375 ;
        RECT 1109.635 104.060 1113.005 104.360 ;
        RECT 1149.180 104.135 1152.480 104.515 ;
        RECT 1153.180 104.135 1156.480 104.515 ;
        RECT 1162.680 104.135 1165.980 104.515 ;
        RECT 1166.680 104.135 1169.980 104.515 ;
        RECT 1101.385 103.325 1101.765 103.705 ;
        RECT 1103.790 103.340 1105.570 103.630 ;
        RECT 1107.045 103.430 1108.235 103.715 ;
        RECT 1111.165 103.310 1112.475 103.630 ;
        RECT 1102.520 102.725 1102.900 103.105 ;
        RECT 1106.265 102.765 1106.645 103.145 ;
        RECT 1108.975 102.755 1109.355 103.135 ;
        RECT 1110.385 102.600 1113.565 102.920 ;
        RECT 1149.180 102.135 1150.465 102.515 ;
        RECT 1168.495 102.135 1169.980 102.515 ;
        RECT 1100.665 101.515 1104.815 101.785 ;
        RECT 1150.685 101.455 1152.205 101.815 ;
        RECT 1100.315 100.010 1104.410 100.015 ;
        RECT 1056.650 100.005 1088.950 100.010 ;
        RECT 1099.195 100.005 1104.410 100.010 ;
        RECT 1002.165 99.990 1006.260 99.995 ;
        RECT 1056.650 99.990 1114.225 100.005 ;
        RECT 1182.295 99.990 1182.675 105.820 ;
        RECT 1191.175 105.770 1195.675 106.080 ;
        RECT 1200.130 105.820 1204.260 106.120 ;
        RECT 1187.135 105.220 1193.525 105.510 ;
        RECT 1186.550 104.640 1197.205 104.975 ;
        RECT 1185.900 104.055 1188.820 104.355 ;
        RECT 1192.365 104.040 1195.735 104.340 ;
        RECT 1184.115 103.305 1184.495 103.685 ;
        RECT 1186.520 103.320 1188.300 103.610 ;
        RECT 1189.775 103.410 1190.965 103.695 ;
        RECT 1193.895 103.290 1195.205 103.610 ;
        RECT 1185.250 102.705 1185.630 103.085 ;
        RECT 1188.995 102.745 1189.375 103.125 ;
        RECT 1191.705 102.735 1192.085 103.115 ;
        RECT 1193.115 102.580 1196.295 102.900 ;
        RECT 1183.045 99.990 1187.140 99.995 ;
        RECT 1197.755 99.990 1198.135 105.820 ;
        RECT 1206.635 105.770 1211.135 106.080 ;
        RECT 1282.820 105.840 1286.950 106.140 ;
        RECT 1289.325 105.790 1293.825 106.100 ;
        RECT 1298.280 105.840 1302.410 106.140 ;
        RECT 1249.320 105.610 1281.065 105.630 ;
        RECT 1202.595 105.220 1208.985 105.510 ;
        RECT 1213.865 105.360 1281.065 105.610 ;
        RECT 1213.865 105.340 1249.775 105.360 ;
        RECT 1285.285 105.240 1291.675 105.530 ;
        RECT 1202.010 104.640 1212.515 104.975 ;
        RECT 1237.485 104.775 1248.035 105.110 ;
        RECT 1276.080 104.795 1280.025 105.130 ;
        RECT 1284.700 104.660 1295.180 104.995 ;
        RECT 1201.360 104.055 1204.280 104.355 ;
        RECT 1207.825 104.040 1211.195 104.340 ;
        RECT 1216.075 104.135 1217.380 104.515 ;
        RECT 1218.080 104.135 1221.380 104.515 ;
        RECT 1222.080 104.135 1225.380 104.515 ;
        RECT 1226.080 104.135 1227.440 104.515 ;
        RECT 1229.415 104.135 1230.880 104.515 ;
        RECT 1231.580 104.135 1234.880 104.515 ;
        RECT 1235.580 104.135 1238.880 104.515 ;
        RECT 1239.580 104.135 1240.760 104.515 ;
        RECT 1254.670 104.155 1255.975 104.535 ;
        RECT 1256.675 104.155 1259.975 104.535 ;
        RECT 1260.675 104.155 1263.975 104.535 ;
        RECT 1264.675 104.155 1266.035 104.535 ;
        RECT 1268.010 104.155 1269.475 104.535 ;
        RECT 1270.175 104.155 1273.475 104.535 ;
        RECT 1274.175 104.155 1277.475 104.535 ;
        RECT 1278.175 104.155 1279.355 104.535 ;
        RECT 1284.050 104.075 1286.970 104.375 ;
        RECT 1290.515 104.060 1293.885 104.360 ;
        RECT 1217.540 103.790 1217.920 103.825 ;
        RECT 1199.575 103.305 1199.955 103.685 ;
        RECT 1201.980 103.320 1203.760 103.610 ;
        RECT 1205.235 103.410 1206.425 103.695 ;
        RECT 1209.355 103.290 1210.665 103.610 ;
        RECT 1217.275 103.480 1220.285 103.790 ;
        RECT 1217.540 103.445 1217.920 103.480 ;
        RECT 1221.540 103.445 1222.630 103.825 ;
        RECT 1225.540 103.820 1225.920 103.825 ;
        RECT 1223.060 103.455 1225.925 103.820 ;
        RECT 1231.040 103.800 1231.420 103.825 ;
        RECT 1231.025 103.480 1233.170 103.800 ;
        RECT 1225.540 103.445 1225.920 103.455 ;
        RECT 1231.040 103.445 1231.420 103.480 ;
        RECT 1234.085 103.445 1235.420 103.825 ;
        RECT 1239.040 103.805 1239.420 103.825 ;
        RECT 1256.135 103.810 1256.515 103.845 ;
        RECT 1236.575 103.485 1239.485 103.805 ;
        RECT 1255.870 103.500 1258.880 103.810 ;
        RECT 1239.040 103.445 1239.420 103.485 ;
        RECT 1256.135 103.465 1256.515 103.500 ;
        RECT 1260.135 103.465 1261.225 103.845 ;
        RECT 1264.135 103.840 1264.515 103.845 ;
        RECT 1261.655 103.475 1264.520 103.840 ;
        RECT 1269.635 103.820 1270.015 103.845 ;
        RECT 1269.620 103.500 1271.765 103.820 ;
        RECT 1264.135 103.465 1264.515 103.475 ;
        RECT 1269.635 103.465 1270.015 103.500 ;
        RECT 1272.680 103.465 1274.015 103.845 ;
        RECT 1277.635 103.825 1278.015 103.845 ;
        RECT 1275.170 103.505 1278.080 103.825 ;
        RECT 1277.635 103.465 1278.015 103.505 ;
        RECT 1282.265 103.325 1282.645 103.705 ;
        RECT 1284.670 103.340 1286.450 103.630 ;
        RECT 1287.925 103.430 1289.115 103.715 ;
        RECT 1292.045 103.310 1293.355 103.630 ;
        RECT 1200.710 102.705 1201.090 103.085 ;
        RECT 1204.455 102.745 1204.835 103.125 ;
        RECT 1207.165 102.735 1207.545 103.115 ;
        RECT 1208.575 102.580 1211.755 102.900 ;
        RECT 1283.400 102.725 1283.780 103.105 ;
        RECT 1287.145 102.765 1287.525 103.145 ;
        RECT 1289.855 102.755 1290.235 103.135 ;
        RECT 1291.265 102.600 1294.445 102.920 ;
        RECT 1215.890 102.135 1217.380 102.515 ;
        RECT 1218.080 102.135 1219.365 102.515 ;
        RECT 1237.395 102.135 1238.880 102.515 ;
        RECT 1239.580 102.135 1240.655 102.515 ;
        RECT 1254.485 102.155 1255.975 102.535 ;
        RECT 1256.675 102.155 1257.960 102.535 ;
        RECT 1275.990 102.155 1277.475 102.535 ;
        RECT 1278.175 102.155 1279.250 102.535 ;
        RECT 1217.540 101.445 1218.630 101.825 ;
        RECT 1219.585 101.455 1221.105 101.815 ;
        RECT 1222.025 101.450 1234.875 101.785 ;
        RECT 1239.040 101.780 1239.420 101.825 ;
        RECT 1238.305 101.480 1239.615 101.780 ;
        RECT 1239.040 101.445 1239.420 101.480 ;
        RECT 1256.135 101.465 1257.225 101.845 ;
        RECT 1258.180 101.475 1259.700 101.835 ;
        RECT 1260.620 101.470 1273.470 101.805 ;
        RECT 1277.635 101.800 1278.015 101.845 ;
        RECT 1276.900 101.500 1278.210 101.800 ;
        RECT 1277.635 101.465 1278.015 101.500 ;
        RECT 1246.695 100.935 1279.645 100.970 ;
        RECT 1214.395 100.605 1279.645 100.935 ;
        RECT 1214.395 100.585 1247.475 100.605 ;
        RECT 1281.440 100.595 1285.700 100.950 ;
        RECT 1279.645 100.010 1285.290 100.015 ;
        RECT 1295.905 100.010 1296.285 105.840 ;
        RECT 1304.785 105.790 1309.285 106.100 ;
        RECT 1300.745 105.240 1307.135 105.530 ;
        RECT 1299.510 104.075 1302.430 104.375 ;
        RECT 1305.975 104.060 1309.345 104.360 ;
        RECT 1297.725 103.325 1298.105 103.705 ;
        RECT 1303.385 103.430 1304.575 103.715 ;
        RECT 1302.605 102.765 1302.985 103.145 ;
        RECT 1306.725 102.600 1309.905 102.920 ;
        RECT 1297.005 101.515 1301.155 101.785 ;
        RECT 1296.655 100.010 1300.750 100.015 ;
        RECT 1252.990 100.005 1285.290 100.010 ;
        RECT 1295.535 100.005 1300.750 100.010 ;
        RECT 1198.505 99.990 1202.600 99.995 ;
        RECT 1252.990 99.990 1310.565 100.005 ;
        RECT 789.245 99.985 794.460 99.990 ;
        RECT 804.705 99.985 809.920 99.990 ;
        RECT 820.165 99.985 917.885 99.990 ;
        RECT 985.585 99.985 990.800 99.990 ;
        RECT 1001.045 99.985 1006.260 99.990 ;
        RECT 1016.505 99.985 1114.225 99.990 ;
        RECT 789.245 99.110 917.885 99.985 ;
        RECT 789.245 99.090 860.415 99.110 ;
        RECT 949.170 99.085 975.825 99.985 ;
        RECT 985.585 99.110 1114.225 99.985 ;
        RECT 985.585 99.090 1056.755 99.110 ;
        RECT 1145.495 99.090 1172.150 99.990 ;
        RECT 1181.925 99.985 1187.140 99.990 ;
        RECT 1197.385 99.985 1202.600 99.990 ;
        RECT 1212.845 99.985 1310.565 99.990 ;
        RECT 1181.925 99.110 1310.565 99.985 ;
        RECT 1181.925 99.090 1253.095 99.110 ;
        RECT 396.530 99.055 467.700 99.075 ;
        RECT 3.635 95.295 76.025 95.320 ;
        RECT 200.000 95.295 272.390 95.320 ;
        RECT -81.535 94.300 -56.100 95.200 ;
        RECT -31.210 94.380 -5.775 95.280 ;
        RECT 3.635 94.420 132.325 95.295 ;
        RECT -79.050 92.120 -77.850 92.500 ;
        RECT -76.095 91.905 -73.820 92.415 ;
        RECT -71.195 91.905 -68.895 92.415 ;
        RECT -66.600 91.905 -64.320 92.415 ;
        RECT -59.525 92.220 -58.290 92.600 ;
        RECT -28.725 92.200 -27.525 92.580 ;
        RECT -25.770 91.985 -23.495 92.495 ;
        RECT -20.870 91.985 -18.570 92.495 ;
        RECT -16.275 91.985 -13.995 92.495 ;
        RECT -9.200 92.300 -7.965 92.680 ;
        RECT -79.050 89.820 -75.790 90.200 ;
        RECT -75.050 89.820 -71.790 90.200 ;
        RECT -65.550 89.820 -62.290 90.200 ;
        RECT -61.550 89.820 -58.290 90.200 ;
        RECT -28.725 89.900 -25.465 90.280 ;
        RECT -24.725 89.900 -21.465 90.280 ;
        RECT -15.225 89.900 -11.965 90.280 ;
        RECT -11.225 89.900 -7.965 90.280 ;
        RECT -78.385 88.235 -56.100 88.245 ;
        RECT -78.385 87.905 -54.560 88.235 ;
        RECT -28.060 87.985 -1.765 88.325 ;
        RECT -56.320 87.885 -54.560 87.905 ;
        RECT 4.005 87.260 4.385 94.420 ;
        RECT 5.835 90.205 9.210 90.605 ;
        RECT 9.580 89.965 9.960 90.345 ;
        RECT 12.295 90.005 12.675 90.385 ;
        RECT 16.480 89.955 16.860 90.335 ;
        RECT 6.905 89.540 8.645 89.830 ;
        RECT 10.695 89.490 11.895 89.780 ;
        RECT 13.405 89.460 16.015 89.885 ;
        RECT 17.615 89.555 17.995 89.935 ;
        RECT 5.150 88.780 18.715 89.095 ;
        RECT 5.145 88.035 18.705 88.335 ;
        RECT 5.165 87.320 11.890 87.620 ;
        RECT 15.590 87.020 18.695 87.295 ;
        RECT 19.465 87.260 19.845 94.420 ;
        RECT 75.970 94.395 132.325 94.420 ;
        RECT 36.105 93.410 73.655 93.435 ;
        RECT 36.105 93.150 101.730 93.410 ;
        RECT 72.955 93.125 101.730 93.150 ;
        RECT 103.400 93.105 110.105 93.405 ;
        RECT 37.615 92.240 39.070 92.620 ;
        RECT 39.810 92.240 41.010 92.620 ;
        RECT 42.765 92.025 45.040 92.535 ;
        RECT 47.665 92.025 49.965 92.535 ;
        RECT 52.260 92.025 54.540 92.535 ;
        RECT 59.335 92.340 60.570 92.720 ;
        RECT 61.310 92.340 62.590 92.720 ;
        RECT 76.260 92.215 77.715 92.595 ;
        RECT 60.750 91.985 61.130 92.020 ;
        RECT 81.410 92.000 83.685 92.510 ;
        RECT 86.310 92.000 88.610 92.510 ;
        RECT 90.905 92.000 93.185 92.510 ;
        RECT 99.955 92.315 101.235 92.695 ;
        RECT 39.250 91.880 39.630 91.920 ;
        RECT 39.180 91.575 42.015 91.880 ;
        RECT 57.995 91.675 61.130 91.985 ;
        RECT 99.395 91.960 99.775 91.995 ;
        RECT 77.895 91.855 78.275 91.895 ;
        RECT 60.750 91.640 61.130 91.675 ;
        RECT 39.250 91.540 39.630 91.575 ;
        RECT 77.825 91.550 80.660 91.855 ;
        RECT 96.640 91.650 99.775 91.960 ;
        RECT 99.395 91.615 99.775 91.650 ;
        RECT 77.895 91.515 78.275 91.550 ;
        RECT 21.295 90.165 24.700 90.605 ;
        RECT 25.040 89.965 25.420 90.345 ;
        RECT 27.755 90.005 28.135 90.385 ;
        RECT 31.940 89.955 32.320 90.335 ;
        RECT 37.775 89.940 39.070 90.320 ;
        RECT 39.810 89.940 43.070 90.320 ;
        RECT 43.810 89.940 47.070 90.320 ;
        RECT 47.810 89.940 48.995 90.320 ;
        RECT 51.260 89.940 52.570 90.320 ;
        RECT 53.310 89.940 56.570 90.320 ;
        RECT 57.310 89.940 60.570 90.320 ;
        RECT 61.310 89.940 62.325 90.320 ;
        RECT 22.365 89.540 24.105 89.830 ;
        RECT 26.155 89.490 27.355 89.780 ;
        RECT 28.865 89.460 31.460 89.835 ;
        RECT 33.075 89.555 33.455 89.935 ;
        RECT 76.420 89.915 77.715 90.295 ;
        RECT 82.455 89.915 85.715 90.295 ;
        RECT 86.455 89.915 87.640 90.295 ;
        RECT 89.905 89.915 91.215 90.295 ;
        RECT 91.955 89.915 95.215 90.295 ;
        RECT 99.955 89.915 100.970 90.295 ;
        RECT 104.035 90.160 107.450 90.580 ;
        RECT 107.780 89.940 108.160 90.320 ;
        RECT 110.495 89.980 110.875 90.360 ;
        RECT 114.680 89.930 115.060 90.310 ;
        RECT 39.250 89.240 39.630 89.620 ;
        RECT 43.250 89.240 43.630 89.620 ;
        RECT 47.250 89.575 47.630 89.620 ;
        RECT 52.750 89.575 53.130 89.620 ;
        RECT 47.200 89.260 53.135 89.575 ;
        RECT 47.250 89.240 47.630 89.260 ;
        RECT 52.750 89.240 53.130 89.260 ;
        RECT 56.750 89.240 57.130 89.620 ;
        RECT 60.750 89.240 61.130 89.620 ;
        RECT 77.895 89.215 78.275 89.595 ;
        RECT 81.895 89.215 82.275 89.595 ;
        RECT 85.895 89.550 86.275 89.595 ;
        RECT 91.395 89.550 91.775 89.595 ;
        RECT 85.845 89.235 91.780 89.550 ;
        RECT 85.895 89.215 86.275 89.235 ;
        RECT 91.395 89.215 91.775 89.235 ;
        RECT 95.395 89.215 95.775 89.595 ;
        RECT 99.395 89.215 99.775 89.595 ;
        RECT 105.105 89.515 106.845 89.805 ;
        RECT 108.895 89.465 110.095 89.755 ;
        RECT 111.605 89.425 114.235 89.880 ;
        RECT 115.815 89.530 116.195 89.910 ;
        RECT 20.605 88.780 34.430 89.080 ;
        RECT 36.105 88.615 52.115 88.990 ;
        RECT 69.985 88.590 90.760 88.965 ;
        RECT 20.610 88.035 39.030 88.335 ;
        RECT 40.475 88.025 67.785 88.365 ;
        RECT 20.090 87.320 27.350 87.620 ;
        RECT 5.145 86.700 9.270 86.970 ;
        RECT 20.645 86.785 24.730 87.055 ;
        RECT 31.050 87.020 34.800 87.295 ;
        RECT 36.105 87.260 62.335 87.650 ;
        RECT 69.015 87.235 100.980 87.625 ;
        RECT 113.790 86.995 116.920 87.270 ;
        RECT 117.665 87.235 118.045 94.395 ;
        RECT 164.960 94.390 190.395 95.290 ;
        RECT 200.000 94.420 328.690 95.295 ;
        RECT 118.905 91.935 125.645 92.235 ;
        RECT 167.445 92.210 168.645 92.590 ;
        RECT 170.400 91.995 172.675 92.505 ;
        RECT 175.300 91.995 177.600 92.505 ;
        RECT 179.895 91.995 182.175 92.505 ;
        RECT 186.970 92.310 188.205 92.690 ;
        RECT 119.495 90.140 122.950 90.580 ;
        RECT 123.240 89.940 123.620 90.320 ;
        RECT 125.955 89.980 126.335 90.360 ;
        RECT 130.140 89.930 130.520 90.310 ;
        RECT 167.445 89.910 170.705 90.290 ;
        RECT 171.445 89.910 174.705 90.290 ;
        RECT 180.945 89.910 184.205 90.290 ;
        RECT 184.945 89.910 188.205 90.290 ;
        RECT 120.565 89.515 122.305 89.805 ;
        RECT 124.355 89.465 125.555 89.755 ;
        RECT 127.065 89.435 129.690 89.845 ;
        RECT 131.275 89.530 131.655 89.910 ;
        RECT 118.310 88.755 134.230 89.055 ;
        RECT 118.845 88.010 135.790 88.310 ;
        RECT 168.110 87.995 194.405 88.335 ;
        RECT 129.250 86.995 136.950 87.270 ;
        RECT 200.370 87.260 200.750 94.420 ;
        RECT 202.200 90.205 205.575 90.605 ;
        RECT 205.945 89.965 206.325 90.345 ;
        RECT 208.660 90.005 209.040 90.385 ;
        RECT 212.845 89.955 213.225 90.335 ;
        RECT 203.270 89.540 205.010 89.830 ;
        RECT 207.060 89.490 208.260 89.780 ;
        RECT 209.770 89.460 212.380 89.885 ;
        RECT 213.980 89.555 214.360 89.935 ;
        RECT 201.515 88.780 215.080 89.095 ;
        RECT 201.510 88.035 215.070 88.335 ;
        RECT 201.530 87.320 208.255 87.620 ;
        RECT 211.955 87.020 215.060 87.295 ;
        RECT 215.830 87.260 216.210 94.420 ;
        RECT 272.335 94.395 328.690 94.420 ;
        RECT 232.470 93.410 270.020 93.435 ;
        RECT 232.470 93.150 298.095 93.410 ;
        RECT 269.320 93.125 298.095 93.150 ;
        RECT 299.765 93.105 306.470 93.405 ;
        RECT 233.980 92.240 235.435 92.620 ;
        RECT 236.175 92.240 237.375 92.620 ;
        RECT 239.130 92.025 241.405 92.535 ;
        RECT 244.030 92.025 246.330 92.535 ;
        RECT 248.625 92.025 250.905 92.535 ;
        RECT 255.700 92.340 256.935 92.720 ;
        RECT 257.675 92.340 258.955 92.720 ;
        RECT 272.625 92.215 274.080 92.595 ;
        RECT 257.115 91.985 257.495 92.020 ;
        RECT 277.775 92.000 280.050 92.510 ;
        RECT 282.675 92.000 284.975 92.510 ;
        RECT 287.270 92.000 289.550 92.510 ;
        RECT 296.320 92.315 297.600 92.695 ;
        RECT 235.615 91.880 235.995 91.920 ;
        RECT 235.545 91.575 238.380 91.880 ;
        RECT 254.360 91.675 257.495 91.985 ;
        RECT 295.760 91.960 296.140 91.995 ;
        RECT 274.260 91.855 274.640 91.895 ;
        RECT 257.115 91.640 257.495 91.675 ;
        RECT 235.615 91.540 235.995 91.575 ;
        RECT 274.190 91.550 277.025 91.855 ;
        RECT 293.005 91.650 296.140 91.960 ;
        RECT 295.760 91.615 296.140 91.650 ;
        RECT 274.260 91.515 274.640 91.550 ;
        RECT 217.660 90.165 221.065 90.605 ;
        RECT 221.405 89.965 221.785 90.345 ;
        RECT 224.120 90.005 224.500 90.385 ;
        RECT 228.305 89.955 228.685 90.335 ;
        RECT 234.140 89.940 235.435 90.320 ;
        RECT 236.175 89.940 239.435 90.320 ;
        RECT 240.175 89.940 243.435 90.320 ;
        RECT 244.175 89.940 245.360 90.320 ;
        RECT 247.625 89.940 248.935 90.320 ;
        RECT 249.675 89.940 252.935 90.320 ;
        RECT 253.675 89.940 256.935 90.320 ;
        RECT 257.675 89.940 258.690 90.320 ;
        RECT 218.730 89.540 220.470 89.830 ;
        RECT 222.520 89.490 223.720 89.780 ;
        RECT 225.230 89.460 227.825 89.835 ;
        RECT 229.440 89.555 229.820 89.935 ;
        RECT 272.785 89.915 274.080 90.295 ;
        RECT 278.820 89.915 282.080 90.295 ;
        RECT 282.820 89.915 284.005 90.295 ;
        RECT 286.270 89.915 287.580 90.295 ;
        RECT 288.320 89.915 291.580 90.295 ;
        RECT 296.320 89.915 297.335 90.295 ;
        RECT 300.400 90.160 303.815 90.580 ;
        RECT 304.145 89.940 304.525 90.320 ;
        RECT 306.860 89.980 307.240 90.360 ;
        RECT 311.045 89.930 311.425 90.310 ;
        RECT 235.615 89.240 235.995 89.620 ;
        RECT 239.615 89.240 239.995 89.620 ;
        RECT 243.615 89.575 243.995 89.620 ;
        RECT 249.115 89.575 249.495 89.620 ;
        RECT 243.565 89.260 249.500 89.575 ;
        RECT 243.615 89.240 243.995 89.260 ;
        RECT 249.115 89.240 249.495 89.260 ;
        RECT 253.115 89.240 253.495 89.620 ;
        RECT 257.115 89.240 257.495 89.620 ;
        RECT 274.260 89.215 274.640 89.595 ;
        RECT 278.260 89.215 278.640 89.595 ;
        RECT 282.260 89.550 282.640 89.595 ;
        RECT 287.760 89.550 288.140 89.595 ;
        RECT 282.210 89.235 288.145 89.550 ;
        RECT 282.260 89.215 282.640 89.235 ;
        RECT 287.760 89.215 288.140 89.235 ;
        RECT 291.760 89.215 292.140 89.595 ;
        RECT 295.760 89.215 296.140 89.595 ;
        RECT 301.470 89.515 303.210 89.805 ;
        RECT 305.260 89.465 306.460 89.755 ;
        RECT 307.970 89.425 310.600 89.880 ;
        RECT 312.180 89.530 312.560 89.910 ;
        RECT 216.970 88.780 230.795 89.080 ;
        RECT 232.470 88.615 248.480 88.990 ;
        RECT 266.350 88.590 287.125 88.965 ;
        RECT 216.975 88.035 235.395 88.335 ;
        RECT 236.840 88.025 264.150 88.365 ;
        RECT 216.455 87.320 223.715 87.620 ;
        RECT 36.105 86.895 54.775 86.905 ;
        RECT 36.105 86.880 66.125 86.895 ;
        RECT 36.105 86.870 93.420 86.880 ;
        RECT 36.105 86.585 102.425 86.870 ;
        RECT 201.510 86.700 205.635 86.970 ;
        RECT 217.010 86.785 221.095 87.055 ;
        RECT 227.415 87.020 231.165 87.295 ;
        RECT 232.470 87.260 258.700 87.650 ;
        RECT 265.380 87.235 297.345 87.625 ;
        RECT 310.155 86.995 313.285 87.270 ;
        RECT 314.030 87.235 314.410 94.395 ;
        RECT 361.350 94.350 386.785 95.250 ;
        RECT 396.400 95.245 468.790 95.270 ;
        RECT 396.400 94.370 525.090 95.245 ;
        RECT 557.670 94.395 583.105 95.295 ;
        RECT 592.775 95.280 665.165 95.305 ;
        RECT 592.775 94.405 721.465 95.280 ;
        RECT 315.270 91.935 322.010 92.235 ;
        RECT 363.835 92.170 365.035 92.550 ;
        RECT 366.790 91.955 369.065 92.465 ;
        RECT 371.690 91.955 373.990 92.465 ;
        RECT 376.285 91.955 378.565 92.465 ;
        RECT 383.360 92.270 384.595 92.650 ;
        RECT 315.860 90.140 319.315 90.580 ;
        RECT 319.605 89.940 319.985 90.320 ;
        RECT 322.320 89.980 322.700 90.360 ;
        RECT 326.505 89.930 326.885 90.310 ;
        RECT 316.930 89.515 318.670 89.805 ;
        RECT 320.720 89.465 321.920 89.755 ;
        RECT 323.430 89.435 326.055 89.845 ;
        RECT 327.640 89.530 328.020 89.910 ;
        RECT 363.835 89.870 367.095 90.250 ;
        RECT 367.835 89.870 371.095 90.250 ;
        RECT 377.335 89.870 380.595 90.250 ;
        RECT 381.335 89.870 384.595 90.250 ;
        RECT 314.675 88.755 330.595 89.055 ;
        RECT 315.210 88.010 332.155 88.310 ;
        RECT 364.500 87.955 390.795 88.295 ;
        RECT 325.615 86.995 333.315 87.270 ;
        RECT 396.770 87.210 397.150 94.370 ;
        RECT 398.600 90.155 401.975 90.555 ;
        RECT 402.345 89.915 402.725 90.295 ;
        RECT 405.060 89.955 405.440 90.335 ;
        RECT 409.245 89.905 409.625 90.285 ;
        RECT 399.670 89.490 401.410 89.780 ;
        RECT 403.460 89.440 404.660 89.730 ;
        RECT 406.170 89.410 408.780 89.835 ;
        RECT 410.380 89.505 410.760 89.885 ;
        RECT 397.915 88.730 411.480 89.045 ;
        RECT 397.910 87.985 411.470 88.285 ;
        RECT 397.930 87.270 404.655 87.570 ;
        RECT 408.355 86.970 411.460 87.245 ;
        RECT 412.230 87.210 412.610 94.370 ;
        RECT 468.735 94.345 525.090 94.370 ;
        RECT 428.870 93.360 466.420 93.385 ;
        RECT 428.870 93.100 494.495 93.360 ;
        RECT 465.720 93.075 494.495 93.100 ;
        RECT 496.165 93.055 502.870 93.355 ;
        RECT 430.380 92.190 431.835 92.570 ;
        RECT 432.575 92.190 433.775 92.570 ;
        RECT 435.530 91.975 437.805 92.485 ;
        RECT 440.430 91.975 442.730 92.485 ;
        RECT 445.025 91.975 447.305 92.485 ;
        RECT 452.100 92.290 453.335 92.670 ;
        RECT 454.075 92.290 455.355 92.670 ;
        RECT 469.025 92.165 470.480 92.545 ;
        RECT 453.515 91.935 453.895 91.970 ;
        RECT 474.175 91.950 476.450 92.460 ;
        RECT 479.075 91.950 481.375 92.460 ;
        RECT 483.670 91.950 485.950 92.460 ;
        RECT 492.720 92.265 494.000 92.645 ;
        RECT 432.015 91.830 432.395 91.870 ;
        RECT 431.945 91.525 434.780 91.830 ;
        RECT 450.760 91.625 453.895 91.935 ;
        RECT 492.160 91.910 492.540 91.945 ;
        RECT 470.660 91.805 471.040 91.845 ;
        RECT 453.515 91.590 453.895 91.625 ;
        RECT 432.015 91.490 432.395 91.525 ;
        RECT 470.590 91.500 473.425 91.805 ;
        RECT 489.405 91.600 492.540 91.910 ;
        RECT 492.160 91.565 492.540 91.600 ;
        RECT 470.660 91.465 471.040 91.500 ;
        RECT 414.060 90.115 417.465 90.555 ;
        RECT 417.805 89.915 418.185 90.295 ;
        RECT 420.520 89.955 420.900 90.335 ;
        RECT 424.705 89.905 425.085 90.285 ;
        RECT 430.540 89.890 431.835 90.270 ;
        RECT 432.575 89.890 435.835 90.270 ;
        RECT 436.575 89.890 439.835 90.270 ;
        RECT 440.575 89.890 441.760 90.270 ;
        RECT 444.025 89.890 445.335 90.270 ;
        RECT 446.075 89.890 449.335 90.270 ;
        RECT 450.075 89.890 453.335 90.270 ;
        RECT 454.075 89.890 455.090 90.270 ;
        RECT 415.130 89.490 416.870 89.780 ;
        RECT 418.920 89.440 420.120 89.730 ;
        RECT 421.630 89.410 424.225 89.785 ;
        RECT 425.840 89.505 426.220 89.885 ;
        RECT 469.185 89.865 470.480 90.245 ;
        RECT 475.220 89.865 478.480 90.245 ;
        RECT 479.220 89.865 480.405 90.245 ;
        RECT 482.670 89.865 483.980 90.245 ;
        RECT 484.720 89.865 487.980 90.245 ;
        RECT 492.720 89.865 493.735 90.245 ;
        RECT 496.800 90.110 500.215 90.530 ;
        RECT 500.545 89.890 500.925 90.270 ;
        RECT 503.260 89.930 503.640 90.310 ;
        RECT 507.445 89.880 507.825 90.260 ;
        RECT 432.015 89.190 432.395 89.570 ;
        RECT 436.015 89.190 436.395 89.570 ;
        RECT 440.015 89.525 440.395 89.570 ;
        RECT 445.515 89.525 445.895 89.570 ;
        RECT 439.965 89.210 445.900 89.525 ;
        RECT 440.015 89.190 440.395 89.210 ;
        RECT 445.515 89.190 445.895 89.210 ;
        RECT 449.515 89.190 449.895 89.570 ;
        RECT 453.515 89.190 453.895 89.570 ;
        RECT 470.660 89.165 471.040 89.545 ;
        RECT 474.660 89.165 475.040 89.545 ;
        RECT 478.660 89.500 479.040 89.545 ;
        RECT 484.160 89.500 484.540 89.545 ;
        RECT 478.610 89.185 484.545 89.500 ;
        RECT 478.660 89.165 479.040 89.185 ;
        RECT 484.160 89.165 484.540 89.185 ;
        RECT 488.160 89.165 488.540 89.545 ;
        RECT 492.160 89.165 492.540 89.545 ;
        RECT 497.870 89.465 499.610 89.755 ;
        RECT 501.660 89.415 502.860 89.705 ;
        RECT 504.370 89.375 507.000 89.830 ;
        RECT 508.580 89.480 508.960 89.860 ;
        RECT 413.370 88.730 427.195 89.030 ;
        RECT 428.870 88.565 444.880 88.940 ;
        RECT 462.750 88.540 483.525 88.915 ;
        RECT 413.375 87.985 431.795 88.285 ;
        RECT 433.240 87.975 460.550 88.315 ;
        RECT 412.855 87.270 420.115 87.570 ;
        RECT 232.470 86.895 251.140 86.905 ;
        RECT 232.470 86.880 262.490 86.895 ;
        RECT 232.470 86.870 289.785 86.880 ;
        RECT 232.470 86.585 298.790 86.870 ;
        RECT 397.910 86.650 402.035 86.920 ;
        RECT 413.410 86.735 417.495 87.005 ;
        RECT 423.815 86.970 427.565 87.245 ;
        RECT 428.870 87.210 455.100 87.600 ;
        RECT 461.780 87.185 493.745 87.575 ;
        RECT 506.555 86.945 509.685 87.220 ;
        RECT 510.430 87.185 510.810 94.345 ;
        RECT 560.155 92.215 561.355 92.595 ;
        RECT 511.670 91.885 518.410 92.185 ;
        RECT 563.110 92.000 565.385 92.510 ;
        RECT 568.010 92.000 570.310 92.510 ;
        RECT 572.605 92.000 574.885 92.510 ;
        RECT 579.680 92.315 580.915 92.695 ;
        RECT 512.260 90.090 515.715 90.530 ;
        RECT 516.005 89.890 516.385 90.270 ;
        RECT 518.720 89.930 519.100 90.310 ;
        RECT 522.905 89.880 523.285 90.260 ;
        RECT 560.155 89.915 563.415 90.295 ;
        RECT 564.155 89.915 567.415 90.295 ;
        RECT 573.655 89.915 576.915 90.295 ;
        RECT 577.655 89.915 580.915 90.295 ;
        RECT 513.330 89.465 515.070 89.755 ;
        RECT 517.120 89.415 518.320 89.705 ;
        RECT 519.830 89.385 522.455 89.795 ;
        RECT 524.040 89.480 524.420 89.860 ;
        RECT 511.075 88.705 526.995 89.005 ;
        RECT 511.610 87.960 528.555 88.260 ;
        RECT 560.820 88.000 587.115 88.340 ;
        RECT 593.145 87.245 593.525 94.405 ;
        RECT 594.975 90.190 598.350 90.590 ;
        RECT 598.720 89.950 599.100 90.330 ;
        RECT 601.435 89.990 601.815 90.370 ;
        RECT 605.620 89.940 606.000 90.320 ;
        RECT 596.045 89.525 597.785 89.815 ;
        RECT 599.835 89.475 601.035 89.765 ;
        RECT 602.545 89.445 605.155 89.870 ;
        RECT 606.755 89.540 607.135 89.920 ;
        RECT 594.290 88.765 607.855 89.080 ;
        RECT 594.285 88.020 607.845 88.320 ;
        RECT 594.305 87.305 601.030 87.605 ;
        RECT 522.015 86.945 529.715 87.220 ;
        RECT 604.730 87.005 607.835 87.280 ;
        RECT 608.605 87.245 608.985 94.405 ;
        RECT 665.110 94.380 721.465 94.405 ;
        RECT 754.035 94.400 779.470 95.300 ;
        RECT 789.115 95.280 861.505 95.305 ;
        RECT 789.115 94.405 917.805 95.280 ;
        RECT 625.245 93.395 662.795 93.420 ;
        RECT 625.245 93.135 690.870 93.395 ;
        RECT 662.095 93.110 690.870 93.135 ;
        RECT 692.540 93.090 699.245 93.390 ;
        RECT 626.755 92.225 628.210 92.605 ;
        RECT 628.950 92.225 630.150 92.605 ;
        RECT 631.905 92.010 634.180 92.520 ;
        RECT 636.805 92.010 639.105 92.520 ;
        RECT 641.400 92.010 643.680 92.520 ;
        RECT 648.475 92.325 649.710 92.705 ;
        RECT 650.450 92.325 651.730 92.705 ;
        RECT 665.400 92.200 666.855 92.580 ;
        RECT 649.890 91.970 650.270 92.005 ;
        RECT 670.550 91.985 672.825 92.495 ;
        RECT 675.450 91.985 677.750 92.495 ;
        RECT 680.045 91.985 682.325 92.495 ;
        RECT 689.095 92.300 690.375 92.680 ;
        RECT 628.390 91.865 628.770 91.905 ;
        RECT 628.320 91.560 631.155 91.865 ;
        RECT 647.135 91.660 650.270 91.970 ;
        RECT 688.535 91.945 688.915 91.980 ;
        RECT 667.035 91.840 667.415 91.880 ;
        RECT 649.890 91.625 650.270 91.660 ;
        RECT 628.390 91.525 628.770 91.560 ;
        RECT 666.965 91.535 669.800 91.840 ;
        RECT 685.780 91.635 688.915 91.945 ;
        RECT 688.535 91.600 688.915 91.635 ;
        RECT 667.035 91.500 667.415 91.535 ;
        RECT 610.435 90.150 613.840 90.590 ;
        RECT 614.180 89.950 614.560 90.330 ;
        RECT 616.895 89.990 617.275 90.370 ;
        RECT 621.080 89.940 621.460 90.320 ;
        RECT 626.915 89.925 628.210 90.305 ;
        RECT 628.950 89.925 632.210 90.305 ;
        RECT 632.950 89.925 636.210 90.305 ;
        RECT 636.950 89.925 638.135 90.305 ;
        RECT 640.400 89.925 641.710 90.305 ;
        RECT 642.450 89.925 645.710 90.305 ;
        RECT 646.450 89.925 649.710 90.305 ;
        RECT 650.450 89.925 651.465 90.305 ;
        RECT 611.505 89.525 613.245 89.815 ;
        RECT 615.295 89.475 616.495 89.765 ;
        RECT 618.005 89.445 620.600 89.820 ;
        RECT 622.215 89.540 622.595 89.920 ;
        RECT 665.560 89.900 666.855 90.280 ;
        RECT 671.595 89.900 674.855 90.280 ;
        RECT 675.595 89.900 676.780 90.280 ;
        RECT 679.045 89.900 680.355 90.280 ;
        RECT 681.095 89.900 684.355 90.280 ;
        RECT 689.095 89.900 690.110 90.280 ;
        RECT 693.175 90.145 696.590 90.565 ;
        RECT 696.920 89.925 697.300 90.305 ;
        RECT 699.635 89.965 700.015 90.345 ;
        RECT 703.820 89.915 704.200 90.295 ;
        RECT 628.390 89.225 628.770 89.605 ;
        RECT 632.390 89.225 632.770 89.605 ;
        RECT 636.390 89.560 636.770 89.605 ;
        RECT 641.890 89.560 642.270 89.605 ;
        RECT 636.340 89.245 642.275 89.560 ;
        RECT 636.390 89.225 636.770 89.245 ;
        RECT 641.890 89.225 642.270 89.245 ;
        RECT 645.890 89.225 646.270 89.605 ;
        RECT 649.890 89.225 650.270 89.605 ;
        RECT 667.035 89.200 667.415 89.580 ;
        RECT 671.035 89.200 671.415 89.580 ;
        RECT 675.035 89.535 675.415 89.580 ;
        RECT 680.535 89.535 680.915 89.580 ;
        RECT 674.985 89.220 680.920 89.535 ;
        RECT 675.035 89.200 675.415 89.220 ;
        RECT 680.535 89.200 680.915 89.220 ;
        RECT 684.535 89.200 684.915 89.580 ;
        RECT 688.535 89.200 688.915 89.580 ;
        RECT 694.245 89.500 695.985 89.790 ;
        RECT 698.035 89.450 699.235 89.740 ;
        RECT 700.745 89.410 703.375 89.865 ;
        RECT 704.955 89.515 705.335 89.895 ;
        RECT 609.745 88.765 623.570 89.065 ;
        RECT 625.245 88.600 641.255 88.975 ;
        RECT 659.125 88.575 679.900 88.950 ;
        RECT 609.750 88.020 628.170 88.320 ;
        RECT 629.615 88.010 656.925 88.350 ;
        RECT 609.230 87.305 616.490 87.605 ;
        RECT 428.870 86.845 447.540 86.855 ;
        RECT 428.870 86.830 458.890 86.845 ;
        RECT 428.870 86.820 486.185 86.830 ;
        RECT 65.860 86.560 102.425 86.585 ;
        RECT 262.225 86.560 298.790 86.585 ;
        RECT 428.870 86.535 495.190 86.820 ;
        RECT 594.285 86.685 598.410 86.955 ;
        RECT 609.785 86.770 613.870 87.040 ;
        RECT 620.190 87.005 623.940 87.280 ;
        RECT 625.245 87.245 651.475 87.635 ;
        RECT 658.155 87.220 690.120 87.610 ;
        RECT 702.930 86.980 706.060 87.255 ;
        RECT 706.805 87.220 707.185 94.380 ;
        RECT 756.520 92.220 757.720 92.600 ;
        RECT 708.045 91.920 714.785 92.220 ;
        RECT 759.475 92.005 761.750 92.515 ;
        RECT 764.375 92.005 766.675 92.515 ;
        RECT 768.970 92.005 771.250 92.515 ;
        RECT 776.045 92.320 777.280 92.700 ;
        RECT 708.635 90.125 712.090 90.565 ;
        RECT 712.380 89.925 712.760 90.305 ;
        RECT 715.095 89.965 715.475 90.345 ;
        RECT 719.280 89.915 719.660 90.295 ;
        RECT 756.520 89.920 759.780 90.300 ;
        RECT 760.520 89.920 763.780 90.300 ;
        RECT 770.020 89.920 773.280 90.300 ;
        RECT 774.020 89.920 777.280 90.300 ;
        RECT 709.705 89.500 711.445 89.790 ;
        RECT 713.495 89.450 714.695 89.740 ;
        RECT 716.205 89.420 718.830 89.830 ;
        RECT 720.415 89.515 720.795 89.895 ;
        RECT 707.450 88.740 723.370 89.040 ;
        RECT 707.985 87.995 724.930 88.295 ;
        RECT 757.185 88.005 783.480 88.345 ;
        RECT 718.390 86.980 726.090 87.255 ;
        RECT 789.485 87.245 789.865 94.405 ;
        RECT 791.315 90.190 794.690 90.590 ;
        RECT 795.060 89.950 795.440 90.330 ;
        RECT 797.775 89.990 798.155 90.370 ;
        RECT 801.960 89.940 802.340 90.320 ;
        RECT 792.385 89.525 794.125 89.815 ;
        RECT 796.175 89.475 797.375 89.765 ;
        RECT 798.885 89.445 801.495 89.870 ;
        RECT 803.095 89.540 803.475 89.920 ;
        RECT 790.630 88.765 804.195 89.080 ;
        RECT 790.625 88.020 804.185 88.320 ;
        RECT 790.645 87.305 797.370 87.605 ;
        RECT 801.070 87.005 804.175 87.280 ;
        RECT 804.945 87.245 805.325 94.405 ;
        RECT 861.450 94.380 917.805 94.405 ;
        RECT 950.420 94.385 975.855 95.285 ;
        RECT 985.455 95.280 1057.845 95.305 ;
        RECT 985.455 94.405 1114.145 95.280 ;
        RECT 821.585 93.395 859.135 93.420 ;
        RECT 821.585 93.135 887.210 93.395 ;
        RECT 858.435 93.110 887.210 93.135 ;
        RECT 888.880 93.090 895.585 93.390 ;
        RECT 823.095 92.225 824.550 92.605 ;
        RECT 825.290 92.225 826.490 92.605 ;
        RECT 828.245 92.010 830.520 92.520 ;
        RECT 833.145 92.010 835.445 92.520 ;
        RECT 837.740 92.010 840.020 92.520 ;
        RECT 844.815 92.325 846.050 92.705 ;
        RECT 846.790 92.325 848.070 92.705 ;
        RECT 861.740 92.200 863.195 92.580 ;
        RECT 846.230 91.970 846.610 92.005 ;
        RECT 866.890 91.985 869.165 92.495 ;
        RECT 871.790 91.985 874.090 92.495 ;
        RECT 876.385 91.985 878.665 92.495 ;
        RECT 885.435 92.300 886.715 92.680 ;
        RECT 824.730 91.865 825.110 91.905 ;
        RECT 824.660 91.560 827.495 91.865 ;
        RECT 843.475 91.660 846.610 91.970 ;
        RECT 884.875 91.945 885.255 91.980 ;
        RECT 863.375 91.840 863.755 91.880 ;
        RECT 846.230 91.625 846.610 91.660 ;
        RECT 824.730 91.525 825.110 91.560 ;
        RECT 863.305 91.535 866.140 91.840 ;
        RECT 882.120 91.635 885.255 91.945 ;
        RECT 884.875 91.600 885.255 91.635 ;
        RECT 863.375 91.500 863.755 91.535 ;
        RECT 806.775 90.150 810.180 90.590 ;
        RECT 810.520 89.950 810.900 90.330 ;
        RECT 813.235 89.990 813.615 90.370 ;
        RECT 817.420 89.940 817.800 90.320 ;
        RECT 823.255 89.925 824.550 90.305 ;
        RECT 825.290 89.925 828.550 90.305 ;
        RECT 829.290 89.925 832.550 90.305 ;
        RECT 833.290 89.925 834.475 90.305 ;
        RECT 836.740 89.925 838.050 90.305 ;
        RECT 838.790 89.925 842.050 90.305 ;
        RECT 842.790 89.925 846.050 90.305 ;
        RECT 846.790 89.925 847.805 90.305 ;
        RECT 807.845 89.525 809.585 89.815 ;
        RECT 811.635 89.475 812.835 89.765 ;
        RECT 814.345 89.445 816.940 89.820 ;
        RECT 818.555 89.540 818.935 89.920 ;
        RECT 861.900 89.900 863.195 90.280 ;
        RECT 867.935 89.900 871.195 90.280 ;
        RECT 871.935 89.900 873.120 90.280 ;
        RECT 875.385 89.900 876.695 90.280 ;
        RECT 877.435 89.900 880.695 90.280 ;
        RECT 885.435 89.900 886.450 90.280 ;
        RECT 889.515 90.145 892.930 90.565 ;
        RECT 893.260 89.925 893.640 90.305 ;
        RECT 895.975 89.965 896.355 90.345 ;
        RECT 900.160 89.915 900.540 90.295 ;
        RECT 824.730 89.225 825.110 89.605 ;
        RECT 828.730 89.225 829.110 89.605 ;
        RECT 832.730 89.560 833.110 89.605 ;
        RECT 838.230 89.560 838.610 89.605 ;
        RECT 832.680 89.245 838.615 89.560 ;
        RECT 832.730 89.225 833.110 89.245 ;
        RECT 838.230 89.225 838.610 89.245 ;
        RECT 842.230 89.225 842.610 89.605 ;
        RECT 846.230 89.225 846.610 89.605 ;
        RECT 863.375 89.200 863.755 89.580 ;
        RECT 867.375 89.200 867.755 89.580 ;
        RECT 871.375 89.535 871.755 89.580 ;
        RECT 876.875 89.535 877.255 89.580 ;
        RECT 871.325 89.220 877.260 89.535 ;
        RECT 871.375 89.200 871.755 89.220 ;
        RECT 876.875 89.200 877.255 89.220 ;
        RECT 880.875 89.200 881.255 89.580 ;
        RECT 884.875 89.200 885.255 89.580 ;
        RECT 890.585 89.500 892.325 89.790 ;
        RECT 894.375 89.450 895.575 89.740 ;
        RECT 897.085 89.410 899.715 89.865 ;
        RECT 901.295 89.515 901.675 89.895 ;
        RECT 806.085 88.765 819.910 89.065 ;
        RECT 821.585 88.600 837.595 88.975 ;
        RECT 855.465 88.575 876.240 88.950 ;
        RECT 806.090 88.020 824.510 88.320 ;
        RECT 825.955 88.010 853.265 88.350 ;
        RECT 805.570 87.305 812.830 87.605 ;
        RECT 625.245 86.880 643.915 86.890 ;
        RECT 625.245 86.865 655.265 86.880 ;
        RECT 625.245 86.855 682.560 86.865 ;
        RECT 625.245 86.570 691.565 86.855 ;
        RECT 790.625 86.685 794.750 86.955 ;
        RECT 806.125 86.770 810.210 87.040 ;
        RECT 816.530 87.005 820.280 87.280 ;
        RECT 821.585 87.245 847.815 87.635 ;
        RECT 854.495 87.220 886.460 87.610 ;
        RECT 899.270 86.980 902.400 87.255 ;
        RECT 903.145 87.220 903.525 94.380 ;
        RECT 904.385 91.920 911.125 92.220 ;
        RECT 952.905 92.205 954.105 92.585 ;
        RECT 955.860 91.990 958.135 92.500 ;
        RECT 960.760 91.990 963.060 92.500 ;
        RECT 965.355 91.990 967.635 92.500 ;
        RECT 972.430 92.305 973.665 92.685 ;
        RECT 904.975 90.125 908.430 90.565 ;
        RECT 908.720 89.925 909.100 90.305 ;
        RECT 911.435 89.965 911.815 90.345 ;
        RECT 915.620 89.915 916.000 90.295 ;
        RECT 952.905 89.905 956.165 90.285 ;
        RECT 956.905 89.905 960.165 90.285 ;
        RECT 966.405 89.905 969.665 90.285 ;
        RECT 970.405 89.905 973.665 90.285 ;
        RECT 906.045 89.500 907.785 89.790 ;
        RECT 909.835 89.450 911.035 89.740 ;
        RECT 912.545 89.420 915.170 89.830 ;
        RECT 916.755 89.515 917.135 89.895 ;
        RECT 903.790 88.740 919.710 89.040 ;
        RECT 904.325 87.995 921.270 88.295 ;
        RECT 953.570 87.990 979.865 88.330 ;
        RECT 914.730 86.980 922.430 87.255 ;
        RECT 985.825 87.245 986.205 94.405 ;
        RECT 987.655 90.190 991.030 90.590 ;
        RECT 991.400 89.950 991.780 90.330 ;
        RECT 994.115 89.990 994.495 90.370 ;
        RECT 998.300 89.940 998.680 90.320 ;
        RECT 988.725 89.525 990.465 89.815 ;
        RECT 992.515 89.475 993.715 89.765 ;
        RECT 995.225 89.445 997.835 89.870 ;
        RECT 999.435 89.540 999.815 89.920 ;
        RECT 986.970 88.765 1000.535 89.080 ;
        RECT 986.965 88.020 1000.525 88.320 ;
        RECT 986.985 87.305 993.710 87.605 ;
        RECT 997.410 87.005 1000.515 87.280 ;
        RECT 1001.285 87.245 1001.665 94.405 ;
        RECT 1057.790 94.380 1114.145 94.405 ;
        RECT 1146.745 94.390 1172.180 95.290 ;
        RECT 1181.795 95.280 1254.185 95.305 ;
        RECT 1181.795 94.405 1310.485 95.280 ;
        RECT 1017.925 93.395 1055.475 93.420 ;
        RECT 1017.925 93.135 1083.550 93.395 ;
        RECT 1054.775 93.110 1083.550 93.135 ;
        RECT 1085.220 93.090 1091.925 93.390 ;
        RECT 1019.435 92.225 1020.890 92.605 ;
        RECT 1021.630 92.225 1022.830 92.605 ;
        RECT 1024.585 92.010 1026.860 92.520 ;
        RECT 1029.485 92.010 1031.785 92.520 ;
        RECT 1034.080 92.010 1036.360 92.520 ;
        RECT 1041.155 92.325 1042.390 92.705 ;
        RECT 1043.130 92.325 1044.410 92.705 ;
        RECT 1058.080 92.200 1059.535 92.580 ;
        RECT 1042.570 91.970 1042.950 92.005 ;
        RECT 1063.230 91.985 1065.505 92.495 ;
        RECT 1068.130 91.985 1070.430 92.495 ;
        RECT 1072.725 91.985 1075.005 92.495 ;
        RECT 1081.775 92.300 1083.055 92.680 ;
        RECT 1021.070 91.865 1021.450 91.905 ;
        RECT 1021.000 91.560 1023.835 91.865 ;
        RECT 1039.815 91.660 1042.950 91.970 ;
        RECT 1081.215 91.945 1081.595 91.980 ;
        RECT 1059.715 91.840 1060.095 91.880 ;
        RECT 1042.570 91.625 1042.950 91.660 ;
        RECT 1021.070 91.525 1021.450 91.560 ;
        RECT 1059.645 91.535 1062.480 91.840 ;
        RECT 1078.460 91.635 1081.595 91.945 ;
        RECT 1081.215 91.600 1081.595 91.635 ;
        RECT 1059.715 91.500 1060.095 91.535 ;
        RECT 1003.115 90.150 1006.520 90.590 ;
        RECT 1006.860 89.950 1007.240 90.330 ;
        RECT 1009.575 89.990 1009.955 90.370 ;
        RECT 1013.760 89.940 1014.140 90.320 ;
        RECT 1019.595 89.925 1020.890 90.305 ;
        RECT 1021.630 89.925 1024.890 90.305 ;
        RECT 1025.630 89.925 1028.890 90.305 ;
        RECT 1029.630 89.925 1030.815 90.305 ;
        RECT 1033.080 89.925 1034.390 90.305 ;
        RECT 1035.130 89.925 1038.390 90.305 ;
        RECT 1039.130 89.925 1042.390 90.305 ;
        RECT 1043.130 89.925 1044.145 90.305 ;
        RECT 1004.185 89.525 1005.925 89.815 ;
        RECT 1007.975 89.475 1009.175 89.765 ;
        RECT 1010.685 89.445 1013.280 89.820 ;
        RECT 1014.895 89.540 1015.275 89.920 ;
        RECT 1058.240 89.900 1059.535 90.280 ;
        RECT 1064.275 89.900 1067.535 90.280 ;
        RECT 1068.275 89.900 1069.460 90.280 ;
        RECT 1071.725 89.900 1073.035 90.280 ;
        RECT 1073.775 89.900 1077.035 90.280 ;
        RECT 1081.775 89.900 1082.790 90.280 ;
        RECT 1085.855 90.145 1089.270 90.565 ;
        RECT 1089.600 89.925 1089.980 90.305 ;
        RECT 1092.315 89.965 1092.695 90.345 ;
        RECT 1096.500 89.915 1096.880 90.295 ;
        RECT 1021.070 89.225 1021.450 89.605 ;
        RECT 1025.070 89.225 1025.450 89.605 ;
        RECT 1029.070 89.560 1029.450 89.605 ;
        RECT 1034.570 89.560 1034.950 89.605 ;
        RECT 1029.020 89.245 1034.955 89.560 ;
        RECT 1029.070 89.225 1029.450 89.245 ;
        RECT 1034.570 89.225 1034.950 89.245 ;
        RECT 1038.570 89.225 1038.950 89.605 ;
        RECT 1042.570 89.225 1042.950 89.605 ;
        RECT 1059.715 89.200 1060.095 89.580 ;
        RECT 1063.715 89.200 1064.095 89.580 ;
        RECT 1067.715 89.535 1068.095 89.580 ;
        RECT 1073.215 89.535 1073.595 89.580 ;
        RECT 1067.665 89.220 1073.600 89.535 ;
        RECT 1067.715 89.200 1068.095 89.220 ;
        RECT 1073.215 89.200 1073.595 89.220 ;
        RECT 1077.215 89.200 1077.595 89.580 ;
        RECT 1081.215 89.200 1081.595 89.580 ;
        RECT 1086.925 89.500 1088.665 89.790 ;
        RECT 1090.715 89.450 1091.915 89.740 ;
        RECT 1093.425 89.410 1096.055 89.865 ;
        RECT 1097.635 89.515 1098.015 89.895 ;
        RECT 1002.425 88.765 1016.250 89.065 ;
        RECT 1017.925 88.600 1033.935 88.975 ;
        RECT 1051.805 88.575 1072.580 88.950 ;
        RECT 1002.430 88.020 1020.850 88.320 ;
        RECT 1022.295 88.010 1049.605 88.350 ;
        RECT 1001.910 87.305 1009.170 87.605 ;
        RECT 821.585 86.880 840.255 86.890 ;
        RECT 821.585 86.865 851.605 86.880 ;
        RECT 821.585 86.855 878.900 86.865 ;
        RECT 821.585 86.570 887.905 86.855 ;
        RECT 986.965 86.685 991.090 86.955 ;
        RECT 1002.465 86.770 1006.550 87.040 ;
        RECT 1012.870 87.005 1016.620 87.280 ;
        RECT 1017.925 87.245 1044.155 87.635 ;
        RECT 1050.835 87.220 1082.800 87.610 ;
        RECT 1095.610 86.980 1098.740 87.255 ;
        RECT 1099.485 87.220 1099.865 94.380 ;
        RECT 1100.725 91.920 1107.465 92.220 ;
        RECT 1149.230 92.210 1150.430 92.590 ;
        RECT 1152.185 91.995 1154.460 92.505 ;
        RECT 1157.085 91.995 1159.385 92.505 ;
        RECT 1161.680 91.995 1163.960 92.505 ;
        RECT 1168.755 92.310 1169.990 92.690 ;
        RECT 1101.315 90.125 1104.770 90.565 ;
        RECT 1105.060 89.925 1105.440 90.305 ;
        RECT 1107.775 89.965 1108.155 90.345 ;
        RECT 1111.960 89.915 1112.340 90.295 ;
        RECT 1149.230 89.910 1152.490 90.290 ;
        RECT 1153.230 89.910 1156.490 90.290 ;
        RECT 1162.730 89.910 1165.990 90.290 ;
        RECT 1166.730 89.910 1169.990 90.290 ;
        RECT 1102.385 89.500 1104.125 89.790 ;
        RECT 1106.175 89.450 1107.375 89.740 ;
        RECT 1108.885 89.420 1111.510 89.830 ;
        RECT 1113.095 89.515 1113.475 89.895 ;
        RECT 1100.130 88.740 1116.050 89.040 ;
        RECT 1100.665 87.995 1117.610 88.295 ;
        RECT 1149.895 87.995 1176.190 88.335 ;
        RECT 1111.070 86.980 1118.770 87.255 ;
        RECT 1182.165 87.245 1182.545 94.405 ;
        RECT 1183.995 90.190 1187.370 90.590 ;
        RECT 1187.740 89.950 1188.120 90.330 ;
        RECT 1190.455 89.990 1190.835 90.370 ;
        RECT 1194.640 89.940 1195.020 90.320 ;
        RECT 1185.065 89.525 1186.805 89.815 ;
        RECT 1188.855 89.475 1190.055 89.765 ;
        RECT 1191.565 89.445 1194.175 89.870 ;
        RECT 1195.775 89.540 1196.155 89.920 ;
        RECT 1183.310 88.765 1196.875 89.080 ;
        RECT 1183.305 88.020 1196.865 88.320 ;
        RECT 1183.325 87.305 1190.050 87.605 ;
        RECT 1193.750 87.005 1196.855 87.280 ;
        RECT 1197.625 87.245 1198.005 94.405 ;
        RECT 1254.130 94.380 1310.485 94.405 ;
        RECT 1214.265 93.395 1251.815 93.420 ;
        RECT 1214.265 93.135 1279.890 93.395 ;
        RECT 1251.115 93.110 1279.890 93.135 ;
        RECT 1281.560 93.090 1288.265 93.390 ;
        RECT 1215.775 92.225 1217.230 92.605 ;
        RECT 1217.970 92.225 1219.170 92.605 ;
        RECT 1220.925 92.010 1223.200 92.520 ;
        RECT 1225.825 92.010 1228.125 92.520 ;
        RECT 1230.420 92.010 1232.700 92.520 ;
        RECT 1237.495 92.325 1238.730 92.705 ;
        RECT 1239.470 92.325 1240.750 92.705 ;
        RECT 1254.420 92.200 1255.875 92.580 ;
        RECT 1256.615 92.200 1257.815 92.580 ;
        RECT 1238.910 91.970 1239.290 92.005 ;
        RECT 1259.570 91.985 1261.845 92.495 ;
        RECT 1264.470 91.985 1266.770 92.495 ;
        RECT 1269.065 91.985 1271.345 92.495 ;
        RECT 1276.140 92.300 1277.375 92.680 ;
        RECT 1278.115 92.300 1279.395 92.680 ;
        RECT 1217.410 91.865 1217.790 91.905 ;
        RECT 1217.340 91.560 1220.175 91.865 ;
        RECT 1236.155 91.660 1239.290 91.970 ;
        RECT 1277.555 91.945 1277.935 91.980 ;
        RECT 1256.055 91.840 1256.435 91.880 ;
        RECT 1238.910 91.625 1239.290 91.660 ;
        RECT 1217.410 91.525 1217.790 91.560 ;
        RECT 1255.985 91.535 1258.820 91.840 ;
        RECT 1274.800 91.635 1277.935 91.945 ;
        RECT 1277.555 91.600 1277.935 91.635 ;
        RECT 1256.055 91.500 1256.435 91.535 ;
        RECT 1199.455 90.150 1202.860 90.590 ;
        RECT 1203.200 89.950 1203.580 90.330 ;
        RECT 1205.915 89.990 1206.295 90.370 ;
        RECT 1210.100 89.940 1210.480 90.320 ;
        RECT 1215.935 89.925 1217.230 90.305 ;
        RECT 1217.970 89.925 1221.230 90.305 ;
        RECT 1221.970 89.925 1225.230 90.305 ;
        RECT 1225.970 89.925 1227.155 90.305 ;
        RECT 1229.420 89.925 1230.730 90.305 ;
        RECT 1231.470 89.925 1234.730 90.305 ;
        RECT 1235.470 89.925 1238.730 90.305 ;
        RECT 1239.470 89.925 1240.485 90.305 ;
        RECT 1200.525 89.525 1202.265 89.815 ;
        RECT 1204.315 89.475 1205.515 89.765 ;
        RECT 1207.025 89.445 1209.620 89.820 ;
        RECT 1211.235 89.540 1211.615 89.920 ;
        RECT 1254.580 89.900 1255.875 90.280 ;
        RECT 1256.615 89.900 1259.875 90.280 ;
        RECT 1260.615 89.900 1263.875 90.280 ;
        RECT 1264.615 89.900 1265.800 90.280 ;
        RECT 1268.065 89.900 1269.375 90.280 ;
        RECT 1270.115 89.900 1273.375 90.280 ;
        RECT 1274.115 89.900 1277.375 90.280 ;
        RECT 1278.115 89.900 1279.130 90.280 ;
        RECT 1282.195 90.145 1285.610 90.565 ;
        RECT 1285.940 89.925 1286.320 90.305 ;
        RECT 1288.655 89.965 1289.035 90.345 ;
        RECT 1292.840 89.915 1293.220 90.295 ;
        RECT 1217.410 89.225 1217.790 89.605 ;
        RECT 1221.410 89.225 1221.790 89.605 ;
        RECT 1225.410 89.560 1225.790 89.605 ;
        RECT 1230.910 89.560 1231.290 89.605 ;
        RECT 1225.360 89.245 1231.295 89.560 ;
        RECT 1225.410 89.225 1225.790 89.245 ;
        RECT 1230.910 89.225 1231.290 89.245 ;
        RECT 1234.910 89.225 1235.290 89.605 ;
        RECT 1238.910 89.225 1239.290 89.605 ;
        RECT 1256.055 89.200 1256.435 89.580 ;
        RECT 1260.055 89.200 1260.435 89.580 ;
        RECT 1264.055 89.535 1264.435 89.580 ;
        RECT 1269.555 89.535 1269.935 89.580 ;
        RECT 1264.005 89.220 1269.940 89.535 ;
        RECT 1264.055 89.200 1264.435 89.220 ;
        RECT 1269.555 89.200 1269.935 89.220 ;
        RECT 1273.555 89.200 1273.935 89.580 ;
        RECT 1277.555 89.200 1277.935 89.580 ;
        RECT 1283.265 89.500 1285.005 89.790 ;
        RECT 1287.055 89.450 1288.255 89.740 ;
        RECT 1289.765 89.410 1292.395 89.865 ;
        RECT 1293.975 89.515 1294.355 89.895 ;
        RECT 1198.765 88.765 1212.590 89.065 ;
        RECT 1214.265 88.600 1230.275 88.975 ;
        RECT 1248.145 88.575 1268.920 88.950 ;
        RECT 1281.545 88.740 1295.160 89.040 ;
        RECT 1198.770 88.020 1217.190 88.320 ;
        RECT 1218.635 88.010 1245.945 88.350 ;
        RECT 1257.280 87.985 1279.835 88.325 ;
        RECT 1280.945 87.995 1295.590 88.295 ;
        RECT 1198.250 87.305 1205.510 87.605 ;
        RECT 1017.925 86.880 1036.595 86.890 ;
        RECT 1017.925 86.865 1047.945 86.880 ;
        RECT 1017.925 86.855 1075.240 86.865 ;
        RECT 1017.925 86.570 1084.245 86.855 ;
        RECT 1183.305 86.685 1187.430 86.955 ;
        RECT 1198.805 86.770 1202.890 87.040 ;
        RECT 1209.210 87.005 1212.960 87.280 ;
        RECT 1214.265 87.245 1240.495 87.635 ;
        RECT 1247.175 87.220 1279.140 87.610 ;
        RECT 1291.950 86.980 1295.080 87.255 ;
        RECT 1295.825 87.220 1296.205 94.380 ;
        RECT 1297.065 91.920 1303.805 92.220 ;
        RECT 1297.655 90.125 1301.110 90.565 ;
        RECT 1304.115 89.965 1304.495 90.345 ;
        RECT 1302.515 89.450 1303.715 89.740 ;
        RECT 1309.435 89.515 1309.815 89.895 ;
        RECT 1296.470 88.740 1312.390 89.040 ;
        RECT 1297.005 87.995 1313.950 88.295 ;
        RECT 1214.265 86.880 1232.935 86.890 ;
        RECT 1214.265 86.865 1244.285 86.880 ;
        RECT 1214.265 86.855 1271.580 86.865 ;
        RECT 1214.265 86.570 1280.585 86.855 ;
        RECT 655.000 86.545 691.565 86.570 ;
        RECT 851.340 86.545 887.905 86.570 ;
        RECT 1047.680 86.545 1084.245 86.570 ;
        RECT 1244.020 86.545 1280.585 86.570 ;
        RECT 458.625 86.510 495.190 86.535 ;
        RECT 6.380 86.125 10.510 86.425 ;
        RECT -59.665 85.285 -56.100 85.295 ;
        RECT -59.665 84.960 -55.305 85.285 ;
        RECT -9.340 85.040 -3.425 85.375 ;
        RECT -6.070 85.020 -3.425 85.040 ;
        RECT -56.260 84.950 -55.305 84.960 ;
        RECT -79.070 84.320 -75.770 84.700 ;
        RECT -75.070 84.320 -71.770 84.700 ;
        RECT -65.570 84.320 -62.270 84.700 ;
        RECT -61.570 84.320 -58.270 84.700 ;
        RECT -28.745 84.400 -25.445 84.780 ;
        RECT -24.745 84.400 -21.445 84.780 ;
        RECT -15.245 84.400 -11.945 84.780 ;
        RECT -11.245 84.400 -7.945 84.780 ;
        RECT -79.070 82.320 -77.785 82.700 ;
        RECT -59.755 82.320 -58.270 82.700 ;
        RECT -28.745 82.400 -27.460 82.780 ;
        RECT -9.430 82.400 -7.945 82.780 ;
        RECT -77.565 81.640 -76.045 82.000 ;
        RECT -27.240 81.720 -25.720 82.080 ;
        RECT 4.005 80.295 4.385 86.125 ;
        RECT 12.885 86.075 17.385 86.385 ;
        RECT 21.840 86.125 25.970 86.425 ;
        RECT 8.845 85.525 15.235 85.815 ;
        RECT 8.260 84.945 18.915 85.280 ;
        RECT 7.610 84.360 10.530 84.660 ;
        RECT 14.075 84.345 17.445 84.645 ;
        RECT 5.825 83.610 6.205 83.990 ;
        RECT 8.230 83.625 10.010 83.915 ;
        RECT 11.485 83.715 12.675 84.000 ;
        RECT 15.605 83.595 16.915 83.915 ;
        RECT 6.960 83.010 7.340 83.390 ;
        RECT 10.705 83.050 11.085 83.430 ;
        RECT 13.415 83.040 13.795 83.420 ;
        RECT 14.825 82.885 18.005 83.205 ;
        RECT 4.755 80.295 8.850 80.300 ;
        RECT 19.465 80.295 19.845 86.125 ;
        RECT 28.345 86.075 32.845 86.385 ;
        RECT 120.040 86.100 124.170 86.400 ;
        RECT 35.575 85.890 71.485 85.915 ;
        RECT 24.305 85.525 30.695 85.815 ;
        RECT 35.575 85.645 102.825 85.890 ;
        RECT 71.080 85.620 102.825 85.645 ;
        RECT 107.045 85.500 113.435 85.790 ;
        RECT 23.720 84.945 34.225 85.280 ;
        RECT 59.195 85.080 69.745 85.415 ;
        RECT 106.460 84.920 116.940 85.255 ;
        RECT 23.070 84.360 25.990 84.660 ;
        RECT 29.535 84.345 32.905 84.645 ;
        RECT 37.785 84.440 39.090 84.820 ;
        RECT 39.790 84.440 43.090 84.820 ;
        RECT 43.790 84.440 47.090 84.820 ;
        RECT 47.790 84.440 49.150 84.820 ;
        RECT 51.125 84.440 52.590 84.820 ;
        RECT 53.290 84.440 56.590 84.820 ;
        RECT 57.290 84.440 60.590 84.820 ;
        RECT 61.290 84.440 62.470 84.820 ;
        RECT 76.430 84.415 77.735 84.795 ;
        RECT 82.435 84.415 85.735 84.795 ;
        RECT 86.435 84.415 87.795 84.795 ;
        RECT 89.770 84.415 91.235 84.795 ;
        RECT 91.935 84.415 95.235 84.795 ;
        RECT 99.935 84.415 101.115 84.795 ;
        RECT 39.250 84.095 39.630 84.130 ;
        RECT 21.285 83.610 21.665 83.990 ;
        RECT 23.690 83.625 25.470 83.915 ;
        RECT 26.945 83.715 28.135 84.000 ;
        RECT 31.065 83.595 32.375 83.915 ;
        RECT 38.985 83.785 41.995 84.095 ;
        RECT 39.250 83.750 39.630 83.785 ;
        RECT 43.250 83.750 44.340 84.130 ;
        RECT 47.250 84.125 47.630 84.130 ;
        RECT 44.770 83.760 47.635 84.125 ;
        RECT 52.750 84.105 53.130 84.130 ;
        RECT 52.735 83.785 54.880 84.105 ;
        RECT 47.250 83.750 47.630 83.760 ;
        RECT 52.750 83.750 53.130 83.785 ;
        RECT 55.795 83.750 57.130 84.130 ;
        RECT 60.750 84.110 61.130 84.130 ;
        RECT 58.285 83.790 61.195 84.110 ;
        RECT 77.895 84.070 78.275 84.105 ;
        RECT 60.750 83.750 61.130 83.790 ;
        RECT 77.630 83.760 80.640 84.070 ;
        RECT 77.895 83.725 78.275 83.760 ;
        RECT 81.895 83.725 82.985 84.105 ;
        RECT 85.895 84.100 86.275 84.105 ;
        RECT 83.415 83.735 86.280 84.100 ;
        RECT 91.395 84.080 91.775 84.105 ;
        RECT 91.380 83.760 93.525 84.080 ;
        RECT 85.895 83.725 86.275 83.735 ;
        RECT 91.395 83.725 91.775 83.760 ;
        RECT 94.440 83.725 95.775 84.105 ;
        RECT 99.395 84.085 99.775 84.105 ;
        RECT 96.930 83.765 99.840 84.085 ;
        RECT 99.395 83.725 99.775 83.765 ;
        RECT 104.025 83.585 104.405 83.965 ;
        RECT 106.430 83.600 108.210 83.890 ;
        RECT 109.685 83.690 110.875 83.975 ;
        RECT 113.805 83.570 115.115 83.890 ;
        RECT 22.420 83.010 22.800 83.390 ;
        RECT 26.165 83.050 26.545 83.430 ;
        RECT 28.875 83.040 29.255 83.420 ;
        RECT 30.285 82.885 33.465 83.205 ;
        RECT 105.160 82.985 105.540 83.365 ;
        RECT 108.905 83.025 109.285 83.405 ;
        RECT 111.615 83.015 111.995 83.395 ;
        RECT 113.025 82.860 116.205 83.180 ;
        RECT 37.600 82.440 39.090 82.820 ;
        RECT 39.790 82.440 41.075 82.820 ;
        RECT 59.105 82.440 60.590 82.820 ;
        RECT 61.290 82.440 62.365 82.820 ;
        RECT 76.245 82.415 77.735 82.795 ;
        RECT 99.935 82.415 101.010 82.795 ;
        RECT 39.250 81.750 40.340 82.130 ;
        RECT 41.295 81.760 42.815 82.120 ;
        RECT 43.735 81.755 56.585 82.090 ;
        RECT 60.750 82.085 61.130 82.130 ;
        RECT 60.015 81.785 61.325 82.085 ;
        RECT 60.750 81.750 61.130 81.785 ;
        RECT 77.895 81.725 78.985 82.105 ;
        RECT 79.940 81.735 81.460 82.095 ;
        RECT 82.380 81.730 95.230 82.065 ;
        RECT 99.395 82.060 99.775 82.105 ;
        RECT 98.660 81.760 99.970 82.060 ;
        RECT 99.395 81.725 99.775 81.760 ;
        RECT 36.105 81.230 69.185 81.240 ;
        RECT 36.105 80.890 101.405 81.230 ;
        RECT 68.455 80.865 101.405 80.890 ;
        RECT 103.200 80.855 107.460 81.210 ;
        RECT 20.215 80.295 24.310 80.300 ;
        RECT 3.635 80.290 8.850 80.295 ;
        RECT 19.095 80.290 24.310 80.295 ;
        RECT 34.555 80.290 74.805 80.295 ;
        RECT 3.635 80.270 74.805 80.290 ;
        RECT 101.405 80.270 107.050 80.275 ;
        RECT 117.665 80.270 118.045 86.100 ;
        RECT 126.545 86.050 131.045 86.360 ;
        RECT 202.745 86.125 206.875 86.425 ;
        RECT 122.505 85.500 128.895 85.790 ;
        RECT 121.920 84.920 137.940 85.255 ;
        RECT 186.830 85.050 192.745 85.385 ;
        RECT 190.100 85.030 192.745 85.050 ;
        RECT 121.270 84.335 124.190 84.635 ;
        RECT 127.735 84.320 131.105 84.620 ;
        RECT 167.425 84.410 170.725 84.790 ;
        RECT 171.425 84.410 174.725 84.790 ;
        RECT 180.925 84.410 184.225 84.790 ;
        RECT 184.925 84.410 188.225 84.790 ;
        RECT 119.485 83.585 119.865 83.965 ;
        RECT 121.890 83.600 123.670 83.890 ;
        RECT 125.145 83.690 126.335 83.975 ;
        RECT 129.265 83.570 130.575 83.890 ;
        RECT 120.620 82.985 121.000 83.365 ;
        RECT 124.365 83.025 124.745 83.405 ;
        RECT 127.075 83.015 127.455 83.395 ;
        RECT 128.485 82.860 131.665 83.180 ;
        RECT 167.425 82.410 168.710 82.790 ;
        RECT 186.740 82.410 188.225 82.790 ;
        RECT 118.765 81.775 122.915 82.045 ;
        RECT 168.930 81.730 170.450 82.090 ;
        RECT 200.370 80.295 200.750 86.125 ;
        RECT 209.250 86.075 213.750 86.385 ;
        RECT 218.205 86.125 222.335 86.425 ;
        RECT 205.210 85.525 211.600 85.815 ;
        RECT 204.625 84.945 215.280 85.280 ;
        RECT 203.975 84.360 206.895 84.660 ;
        RECT 210.440 84.345 213.810 84.645 ;
        RECT 202.190 83.610 202.570 83.990 ;
        RECT 204.595 83.625 206.375 83.915 ;
        RECT 207.850 83.715 209.040 84.000 ;
        RECT 211.970 83.595 213.280 83.915 ;
        RECT 203.325 83.010 203.705 83.390 ;
        RECT 207.070 83.050 207.450 83.430 ;
        RECT 209.780 83.040 210.160 83.420 ;
        RECT 211.190 82.885 214.370 83.205 ;
        RECT 201.120 80.295 205.215 80.300 ;
        RECT 215.830 80.295 216.210 86.125 ;
        RECT 224.710 86.075 229.210 86.385 ;
        RECT 316.405 86.100 320.535 86.400 ;
        RECT 231.940 85.890 267.850 85.915 ;
        RECT 220.670 85.525 227.060 85.815 ;
        RECT 231.940 85.645 299.190 85.890 ;
        RECT 267.445 85.620 299.190 85.645 ;
        RECT 303.410 85.500 309.800 85.790 ;
        RECT 220.085 84.945 230.590 85.280 ;
        RECT 255.560 85.080 266.110 85.415 ;
        RECT 302.825 84.920 313.305 85.255 ;
        RECT 219.435 84.360 222.355 84.660 ;
        RECT 225.900 84.345 229.270 84.645 ;
        RECT 234.150 84.440 235.455 84.820 ;
        RECT 236.155 84.440 239.455 84.820 ;
        RECT 240.155 84.440 243.455 84.820 ;
        RECT 244.155 84.440 245.515 84.820 ;
        RECT 247.490 84.440 248.955 84.820 ;
        RECT 249.655 84.440 252.955 84.820 ;
        RECT 253.655 84.440 256.955 84.820 ;
        RECT 257.655 84.440 258.835 84.820 ;
        RECT 272.795 84.415 274.100 84.795 ;
        RECT 278.800 84.415 282.100 84.795 ;
        RECT 282.800 84.415 284.160 84.795 ;
        RECT 286.135 84.415 287.600 84.795 ;
        RECT 288.300 84.415 291.600 84.795 ;
        RECT 296.300 84.415 297.480 84.795 ;
        RECT 235.615 84.095 235.995 84.130 ;
        RECT 217.650 83.610 218.030 83.990 ;
        RECT 220.055 83.625 221.835 83.915 ;
        RECT 223.310 83.715 224.500 84.000 ;
        RECT 227.430 83.595 228.740 83.915 ;
        RECT 235.350 83.785 238.360 84.095 ;
        RECT 235.615 83.750 235.995 83.785 ;
        RECT 239.615 83.750 240.705 84.130 ;
        RECT 243.615 84.125 243.995 84.130 ;
        RECT 241.135 83.760 244.000 84.125 ;
        RECT 249.115 84.105 249.495 84.130 ;
        RECT 249.100 83.785 251.245 84.105 ;
        RECT 243.615 83.750 243.995 83.760 ;
        RECT 249.115 83.750 249.495 83.785 ;
        RECT 252.160 83.750 253.495 84.130 ;
        RECT 257.115 84.110 257.495 84.130 ;
        RECT 254.650 83.790 257.560 84.110 ;
        RECT 274.260 84.070 274.640 84.105 ;
        RECT 257.115 83.750 257.495 83.790 ;
        RECT 273.995 83.760 277.005 84.070 ;
        RECT 274.260 83.725 274.640 83.760 ;
        RECT 278.260 83.725 279.350 84.105 ;
        RECT 282.260 84.100 282.640 84.105 ;
        RECT 279.780 83.735 282.645 84.100 ;
        RECT 287.760 84.080 288.140 84.105 ;
        RECT 287.745 83.760 289.890 84.080 ;
        RECT 282.260 83.725 282.640 83.735 ;
        RECT 287.760 83.725 288.140 83.760 ;
        RECT 290.805 83.725 292.140 84.105 ;
        RECT 295.760 84.085 296.140 84.105 ;
        RECT 293.295 83.765 296.205 84.085 ;
        RECT 295.760 83.725 296.140 83.765 ;
        RECT 300.390 83.585 300.770 83.965 ;
        RECT 302.795 83.600 304.575 83.890 ;
        RECT 306.050 83.690 307.240 83.975 ;
        RECT 310.170 83.570 311.480 83.890 ;
        RECT 218.785 83.010 219.165 83.390 ;
        RECT 222.530 83.050 222.910 83.430 ;
        RECT 225.240 83.040 225.620 83.420 ;
        RECT 226.650 82.885 229.830 83.205 ;
        RECT 301.525 82.985 301.905 83.365 ;
        RECT 305.270 83.025 305.650 83.405 ;
        RECT 307.980 83.015 308.360 83.395 ;
        RECT 309.390 82.860 312.570 83.180 ;
        RECT 233.965 82.440 235.455 82.820 ;
        RECT 236.155 82.440 237.440 82.820 ;
        RECT 255.470 82.440 256.955 82.820 ;
        RECT 257.655 82.440 258.730 82.820 ;
        RECT 272.610 82.415 274.100 82.795 ;
        RECT 296.300 82.415 297.375 82.795 ;
        RECT 235.615 81.750 236.705 82.130 ;
        RECT 237.660 81.760 239.180 82.120 ;
        RECT 240.100 81.755 252.950 82.090 ;
        RECT 257.115 82.085 257.495 82.130 ;
        RECT 256.380 81.785 257.690 82.085 ;
        RECT 257.115 81.750 257.495 81.785 ;
        RECT 274.260 81.725 275.350 82.105 ;
        RECT 276.305 81.735 277.825 82.095 ;
        RECT 278.745 81.730 291.595 82.065 ;
        RECT 295.760 82.060 296.140 82.105 ;
        RECT 295.025 81.760 296.335 82.060 ;
        RECT 295.760 81.725 296.140 81.760 ;
        RECT 232.470 81.230 265.550 81.240 ;
        RECT 232.470 80.890 297.770 81.230 ;
        RECT 264.820 80.865 297.770 80.890 ;
        RECT 299.565 80.855 303.825 81.210 ;
        RECT 216.580 80.295 220.675 80.300 ;
        RECT 200.000 80.290 205.215 80.295 ;
        RECT 215.460 80.290 220.675 80.295 ;
        RECT 230.920 80.290 271.170 80.295 ;
        RECT 118.415 80.270 122.510 80.275 ;
        RECT 3.635 80.265 107.050 80.270 ;
        RECT 117.295 80.265 122.510 80.270 ;
        RECT 200.000 80.270 271.170 80.290 ;
        RECT 297.770 80.270 303.415 80.275 ;
        RECT 314.030 80.270 314.410 86.100 ;
        RECT 322.910 86.050 327.410 86.360 ;
        RECT 399.145 86.075 403.275 86.375 ;
        RECT 318.870 85.500 325.260 85.790 ;
        RECT 318.285 84.920 334.305 85.255 ;
        RECT 383.220 85.010 389.135 85.345 ;
        RECT 386.490 84.990 389.135 85.010 ;
        RECT 317.635 84.335 320.555 84.635 ;
        RECT 324.100 84.320 327.470 84.620 ;
        RECT 363.815 84.370 367.115 84.750 ;
        RECT 367.815 84.370 371.115 84.750 ;
        RECT 377.315 84.370 380.615 84.750 ;
        RECT 381.315 84.370 384.615 84.750 ;
        RECT 315.850 83.585 316.230 83.965 ;
        RECT 318.255 83.600 320.035 83.890 ;
        RECT 321.510 83.690 322.700 83.975 ;
        RECT 325.630 83.570 326.940 83.890 ;
        RECT 316.985 82.985 317.365 83.365 ;
        RECT 320.730 83.025 321.110 83.405 ;
        RECT 323.440 83.015 323.820 83.395 ;
        RECT 324.850 82.860 328.030 83.180 ;
        RECT 363.815 82.370 365.100 82.750 ;
        RECT 383.130 82.370 384.615 82.750 ;
        RECT 315.130 81.775 319.280 82.045 ;
        RECT 365.320 81.690 366.840 82.050 ;
        RECT 314.780 80.270 318.875 80.275 ;
        RECT 200.000 80.265 303.415 80.270 ;
        RECT 313.660 80.265 318.875 80.270 ;
        RECT -82.755 79.275 -56.100 80.175 ;
        RECT -32.430 79.355 -5.775 80.255 ;
        RECT 3.635 79.395 132.325 80.265 ;
        RECT 74.750 79.370 132.325 79.395 ;
        RECT 163.740 79.365 190.395 80.265 ;
        RECT 200.000 79.395 328.690 80.265 ;
        RECT 396.770 80.245 397.150 86.075 ;
        RECT 405.650 86.025 410.150 86.335 ;
        RECT 414.605 86.075 418.735 86.375 ;
        RECT 401.610 85.475 408.000 85.765 ;
        RECT 401.025 84.895 411.680 85.230 ;
        RECT 400.375 84.310 403.295 84.610 ;
        RECT 406.840 84.295 410.210 84.595 ;
        RECT 398.590 83.560 398.970 83.940 ;
        RECT 400.995 83.575 402.775 83.865 ;
        RECT 404.250 83.665 405.440 83.950 ;
        RECT 408.370 83.545 409.680 83.865 ;
        RECT 399.725 82.960 400.105 83.340 ;
        RECT 403.470 83.000 403.850 83.380 ;
        RECT 406.180 82.990 406.560 83.370 ;
        RECT 407.590 82.835 410.770 83.155 ;
        RECT 397.520 80.245 401.615 80.250 ;
        RECT 412.230 80.245 412.610 86.075 ;
        RECT 421.110 86.025 425.610 86.335 ;
        RECT 512.805 86.050 516.935 86.350 ;
        RECT 428.340 85.840 464.250 85.865 ;
        RECT 417.070 85.475 423.460 85.765 ;
        RECT 428.340 85.595 495.590 85.840 ;
        RECT 463.845 85.570 495.590 85.595 ;
        RECT 499.810 85.450 506.200 85.740 ;
        RECT 416.485 84.895 426.990 85.230 ;
        RECT 451.960 85.030 462.510 85.365 ;
        RECT 499.225 84.870 509.705 85.205 ;
        RECT 415.835 84.310 418.755 84.610 ;
        RECT 422.300 84.295 425.670 84.595 ;
        RECT 430.550 84.390 431.855 84.770 ;
        RECT 432.555 84.390 435.855 84.770 ;
        RECT 436.555 84.390 439.855 84.770 ;
        RECT 440.555 84.390 441.915 84.770 ;
        RECT 443.890 84.390 445.355 84.770 ;
        RECT 446.055 84.390 449.355 84.770 ;
        RECT 450.055 84.390 453.355 84.770 ;
        RECT 454.055 84.390 455.235 84.770 ;
        RECT 469.195 84.365 470.500 84.745 ;
        RECT 475.200 84.365 478.500 84.745 ;
        RECT 479.200 84.365 480.560 84.745 ;
        RECT 482.535 84.365 484.000 84.745 ;
        RECT 484.700 84.365 488.000 84.745 ;
        RECT 492.700 84.365 493.880 84.745 ;
        RECT 432.015 84.045 432.395 84.080 ;
        RECT 414.050 83.560 414.430 83.940 ;
        RECT 416.455 83.575 418.235 83.865 ;
        RECT 419.710 83.665 420.900 83.950 ;
        RECT 423.830 83.545 425.140 83.865 ;
        RECT 431.750 83.735 434.760 84.045 ;
        RECT 432.015 83.700 432.395 83.735 ;
        RECT 436.015 83.700 437.105 84.080 ;
        RECT 440.015 84.075 440.395 84.080 ;
        RECT 437.535 83.710 440.400 84.075 ;
        RECT 445.515 84.055 445.895 84.080 ;
        RECT 445.500 83.735 447.645 84.055 ;
        RECT 440.015 83.700 440.395 83.710 ;
        RECT 445.515 83.700 445.895 83.735 ;
        RECT 448.560 83.700 449.895 84.080 ;
        RECT 453.515 84.060 453.895 84.080 ;
        RECT 451.050 83.740 453.960 84.060 ;
        RECT 470.660 84.020 471.040 84.055 ;
        RECT 453.515 83.700 453.895 83.740 ;
        RECT 470.395 83.710 473.405 84.020 ;
        RECT 470.660 83.675 471.040 83.710 ;
        RECT 474.660 83.675 475.750 84.055 ;
        RECT 478.660 84.050 479.040 84.055 ;
        RECT 476.180 83.685 479.045 84.050 ;
        RECT 484.160 84.030 484.540 84.055 ;
        RECT 484.145 83.710 486.290 84.030 ;
        RECT 478.660 83.675 479.040 83.685 ;
        RECT 484.160 83.675 484.540 83.710 ;
        RECT 487.205 83.675 488.540 84.055 ;
        RECT 492.160 84.035 492.540 84.055 ;
        RECT 489.695 83.715 492.605 84.035 ;
        RECT 492.160 83.675 492.540 83.715 ;
        RECT 496.790 83.535 497.170 83.915 ;
        RECT 499.195 83.550 500.975 83.840 ;
        RECT 502.450 83.640 503.640 83.925 ;
        RECT 506.570 83.520 507.880 83.840 ;
        RECT 415.185 82.960 415.565 83.340 ;
        RECT 418.930 83.000 419.310 83.380 ;
        RECT 421.640 82.990 422.020 83.370 ;
        RECT 423.050 82.835 426.230 83.155 ;
        RECT 497.925 82.935 498.305 83.315 ;
        RECT 501.670 82.975 502.050 83.355 ;
        RECT 504.380 82.965 504.760 83.345 ;
        RECT 505.790 82.810 508.970 83.130 ;
        RECT 430.365 82.390 431.855 82.770 ;
        RECT 432.555 82.390 433.840 82.770 ;
        RECT 451.870 82.390 453.355 82.770 ;
        RECT 454.055 82.390 455.130 82.770 ;
        RECT 469.010 82.365 470.500 82.745 ;
        RECT 492.700 82.365 493.775 82.745 ;
        RECT 432.015 81.700 433.105 82.080 ;
        RECT 434.060 81.710 435.580 82.070 ;
        RECT 436.500 81.705 449.350 82.040 ;
        RECT 453.515 82.035 453.895 82.080 ;
        RECT 452.780 81.735 454.090 82.035 ;
        RECT 453.515 81.700 453.895 81.735 ;
        RECT 470.660 81.675 471.750 82.055 ;
        RECT 472.705 81.685 474.225 82.045 ;
        RECT 475.145 81.680 487.995 82.015 ;
        RECT 492.160 82.010 492.540 82.055 ;
        RECT 491.425 81.710 492.735 82.010 ;
        RECT 492.160 81.675 492.540 81.710 ;
        RECT 428.870 81.180 461.950 81.190 ;
        RECT 428.870 80.840 494.170 81.180 ;
        RECT 461.220 80.815 494.170 80.840 ;
        RECT 495.965 80.805 500.225 81.160 ;
        RECT 412.980 80.245 417.075 80.250 ;
        RECT 396.400 80.240 401.615 80.245 ;
        RECT 411.860 80.240 417.075 80.245 ;
        RECT 427.320 80.240 467.570 80.245 ;
        RECT 271.115 79.370 328.690 79.395 ;
        RECT 360.130 79.325 386.785 80.225 ;
        RECT 396.400 80.220 467.570 80.240 ;
        RECT 494.170 80.220 499.815 80.225 ;
        RECT 510.430 80.220 510.810 86.050 ;
        RECT 519.310 86.000 523.810 86.310 ;
        RECT 595.520 86.110 599.650 86.410 ;
        RECT 515.270 85.450 521.660 85.740 ;
        RECT 514.685 84.870 530.705 85.205 ;
        RECT 579.540 85.055 585.455 85.390 ;
        RECT 582.810 85.035 585.455 85.055 ;
        RECT 514.035 84.285 516.955 84.585 ;
        RECT 520.500 84.270 523.870 84.570 ;
        RECT 560.135 84.415 563.435 84.795 ;
        RECT 564.135 84.415 567.435 84.795 ;
        RECT 573.635 84.415 576.935 84.795 ;
        RECT 577.635 84.415 580.935 84.795 ;
        RECT 512.250 83.535 512.630 83.915 ;
        RECT 514.655 83.550 516.435 83.840 ;
        RECT 517.910 83.640 519.100 83.925 ;
        RECT 522.030 83.520 523.340 83.840 ;
        RECT 513.385 82.935 513.765 83.315 ;
        RECT 517.130 82.975 517.510 83.355 ;
        RECT 519.840 82.965 520.220 83.345 ;
        RECT 521.250 82.810 524.430 83.130 ;
        RECT 560.135 82.415 561.420 82.795 ;
        RECT 579.450 82.415 580.935 82.795 ;
        RECT 511.530 81.725 515.680 81.995 ;
        RECT 561.640 81.735 563.160 82.095 ;
        RECT 593.145 80.280 593.525 86.110 ;
        RECT 602.025 86.060 606.525 86.370 ;
        RECT 610.980 86.110 615.110 86.410 ;
        RECT 597.985 85.510 604.375 85.800 ;
        RECT 597.400 84.930 608.055 85.265 ;
        RECT 596.750 84.345 599.670 84.645 ;
        RECT 603.215 84.330 606.585 84.630 ;
        RECT 594.965 83.595 595.345 83.975 ;
        RECT 597.370 83.610 599.150 83.900 ;
        RECT 600.625 83.700 601.815 83.985 ;
        RECT 604.745 83.580 606.055 83.900 ;
        RECT 596.100 82.995 596.480 83.375 ;
        RECT 599.845 83.035 600.225 83.415 ;
        RECT 602.555 83.025 602.935 83.405 ;
        RECT 603.965 82.870 607.145 83.190 ;
        RECT 593.895 80.280 597.990 80.285 ;
        RECT 608.605 80.280 608.985 86.110 ;
        RECT 617.485 86.060 621.985 86.370 ;
        RECT 709.180 86.085 713.310 86.385 ;
        RECT 624.715 85.875 660.625 85.900 ;
        RECT 613.445 85.510 619.835 85.800 ;
        RECT 624.715 85.630 691.965 85.875 ;
        RECT 660.220 85.605 691.965 85.630 ;
        RECT 696.185 85.485 702.575 85.775 ;
        RECT 612.860 84.930 623.365 85.265 ;
        RECT 648.335 85.065 658.885 85.400 ;
        RECT 695.600 84.905 706.080 85.240 ;
        RECT 612.210 84.345 615.130 84.645 ;
        RECT 618.675 84.330 622.045 84.630 ;
        RECT 626.925 84.425 628.230 84.805 ;
        RECT 628.930 84.425 632.230 84.805 ;
        RECT 632.930 84.425 636.230 84.805 ;
        RECT 636.930 84.425 638.290 84.805 ;
        RECT 640.265 84.425 641.730 84.805 ;
        RECT 642.430 84.425 645.730 84.805 ;
        RECT 646.430 84.425 649.730 84.805 ;
        RECT 650.430 84.425 651.610 84.805 ;
        RECT 665.570 84.400 666.875 84.780 ;
        RECT 671.575 84.400 674.875 84.780 ;
        RECT 675.575 84.400 676.935 84.780 ;
        RECT 678.910 84.400 680.375 84.780 ;
        RECT 681.075 84.400 684.375 84.780 ;
        RECT 689.075 84.400 690.255 84.780 ;
        RECT 628.390 84.080 628.770 84.115 ;
        RECT 610.425 83.595 610.805 83.975 ;
        RECT 612.830 83.610 614.610 83.900 ;
        RECT 616.085 83.700 617.275 83.985 ;
        RECT 620.205 83.580 621.515 83.900 ;
        RECT 628.125 83.770 631.135 84.080 ;
        RECT 628.390 83.735 628.770 83.770 ;
        RECT 632.390 83.735 633.480 84.115 ;
        RECT 636.390 84.110 636.770 84.115 ;
        RECT 633.910 83.745 636.775 84.110 ;
        RECT 641.890 84.090 642.270 84.115 ;
        RECT 641.875 83.770 644.020 84.090 ;
        RECT 636.390 83.735 636.770 83.745 ;
        RECT 641.890 83.735 642.270 83.770 ;
        RECT 644.935 83.735 646.270 84.115 ;
        RECT 649.890 84.095 650.270 84.115 ;
        RECT 647.425 83.775 650.335 84.095 ;
        RECT 667.035 84.055 667.415 84.090 ;
        RECT 649.890 83.735 650.270 83.775 ;
        RECT 666.770 83.745 669.780 84.055 ;
        RECT 667.035 83.710 667.415 83.745 ;
        RECT 671.035 83.710 672.125 84.090 ;
        RECT 675.035 84.085 675.415 84.090 ;
        RECT 672.555 83.720 675.420 84.085 ;
        RECT 680.535 84.065 680.915 84.090 ;
        RECT 680.520 83.745 682.665 84.065 ;
        RECT 675.035 83.710 675.415 83.720 ;
        RECT 680.535 83.710 680.915 83.745 ;
        RECT 683.580 83.710 684.915 84.090 ;
        RECT 688.535 84.070 688.915 84.090 ;
        RECT 686.070 83.750 688.980 84.070 ;
        RECT 688.535 83.710 688.915 83.750 ;
        RECT 693.165 83.570 693.545 83.950 ;
        RECT 695.570 83.585 697.350 83.875 ;
        RECT 698.825 83.675 700.015 83.960 ;
        RECT 702.945 83.555 704.255 83.875 ;
        RECT 611.560 82.995 611.940 83.375 ;
        RECT 615.305 83.035 615.685 83.415 ;
        RECT 618.015 83.025 618.395 83.405 ;
        RECT 619.425 82.870 622.605 83.190 ;
        RECT 694.300 82.970 694.680 83.350 ;
        RECT 698.045 83.010 698.425 83.390 ;
        RECT 700.755 83.000 701.135 83.380 ;
        RECT 702.165 82.845 705.345 83.165 ;
        RECT 626.740 82.425 628.230 82.805 ;
        RECT 628.930 82.425 630.215 82.805 ;
        RECT 648.245 82.425 649.730 82.805 ;
        RECT 650.430 82.425 651.505 82.805 ;
        RECT 665.385 82.400 666.875 82.780 ;
        RECT 689.075 82.400 690.150 82.780 ;
        RECT 628.390 81.735 629.480 82.115 ;
        RECT 630.435 81.745 631.955 82.105 ;
        RECT 632.875 81.740 645.725 82.075 ;
        RECT 649.890 82.070 650.270 82.115 ;
        RECT 649.155 81.770 650.465 82.070 ;
        RECT 649.890 81.735 650.270 81.770 ;
        RECT 667.035 81.710 668.125 82.090 ;
        RECT 669.080 81.720 670.600 82.080 ;
        RECT 671.520 81.715 684.370 82.050 ;
        RECT 688.535 82.045 688.915 82.090 ;
        RECT 687.800 81.745 689.110 82.045 ;
        RECT 688.535 81.710 688.915 81.745 ;
        RECT 625.245 81.215 658.325 81.225 ;
        RECT 625.245 80.875 690.545 81.215 ;
        RECT 657.595 80.850 690.545 80.875 ;
        RECT 692.340 80.840 696.600 81.195 ;
        RECT 609.355 80.280 613.450 80.285 ;
        RECT 592.775 80.275 597.990 80.280 ;
        RECT 608.235 80.275 613.450 80.280 ;
        RECT 623.695 80.275 663.945 80.280 ;
        RECT 511.180 80.220 515.275 80.225 ;
        RECT 396.400 80.215 499.815 80.220 ;
        RECT 510.060 80.215 515.275 80.220 ;
        RECT 396.400 79.345 525.090 80.215 ;
        RECT 556.450 79.370 583.105 80.270 ;
        RECT 592.775 80.255 663.945 80.275 ;
        RECT 690.545 80.255 696.190 80.260 ;
        RECT 706.805 80.255 707.185 86.085 ;
        RECT 715.685 86.035 720.185 86.345 ;
        RECT 791.860 86.110 795.990 86.410 ;
        RECT 711.645 85.485 718.035 85.775 ;
        RECT 711.060 84.905 727.080 85.240 ;
        RECT 775.905 85.060 781.820 85.395 ;
        RECT 779.175 85.040 781.820 85.060 ;
        RECT 710.410 84.320 713.330 84.620 ;
        RECT 716.875 84.305 720.245 84.605 ;
        RECT 756.500 84.420 759.800 84.800 ;
        RECT 760.500 84.420 763.800 84.800 ;
        RECT 770.000 84.420 773.300 84.800 ;
        RECT 774.000 84.420 777.300 84.800 ;
        RECT 708.625 83.570 709.005 83.950 ;
        RECT 711.030 83.585 712.810 83.875 ;
        RECT 714.285 83.675 715.475 83.960 ;
        RECT 718.405 83.555 719.715 83.875 ;
        RECT 709.760 82.970 710.140 83.350 ;
        RECT 713.505 83.010 713.885 83.390 ;
        RECT 716.215 83.000 716.595 83.380 ;
        RECT 717.625 82.845 720.805 83.165 ;
        RECT 756.500 82.420 757.785 82.800 ;
        RECT 775.815 82.420 777.300 82.800 ;
        RECT 707.905 81.760 712.055 82.030 ;
        RECT 758.005 81.740 759.525 82.100 ;
        RECT 789.485 80.280 789.865 86.110 ;
        RECT 798.365 86.060 802.865 86.370 ;
        RECT 807.320 86.110 811.450 86.410 ;
        RECT 794.325 85.510 800.715 85.800 ;
        RECT 793.740 84.930 804.395 85.265 ;
        RECT 793.090 84.345 796.010 84.645 ;
        RECT 799.555 84.330 802.925 84.630 ;
        RECT 791.305 83.595 791.685 83.975 ;
        RECT 793.710 83.610 795.490 83.900 ;
        RECT 796.965 83.700 798.155 83.985 ;
        RECT 801.085 83.580 802.395 83.900 ;
        RECT 792.440 82.995 792.820 83.375 ;
        RECT 796.185 83.035 796.565 83.415 ;
        RECT 798.895 83.025 799.275 83.405 ;
        RECT 800.305 82.870 803.485 83.190 ;
        RECT 790.235 80.280 794.330 80.285 ;
        RECT 804.945 80.280 805.325 86.110 ;
        RECT 813.825 86.060 818.325 86.370 ;
        RECT 905.520 86.085 909.650 86.385 ;
        RECT 821.055 85.875 856.965 85.900 ;
        RECT 809.785 85.510 816.175 85.800 ;
        RECT 821.055 85.630 888.305 85.875 ;
        RECT 856.560 85.605 888.305 85.630 ;
        RECT 892.525 85.485 898.915 85.775 ;
        RECT 809.200 84.930 819.705 85.265 ;
        RECT 844.675 85.065 855.225 85.400 ;
        RECT 891.940 84.905 902.420 85.240 ;
        RECT 808.550 84.345 811.470 84.645 ;
        RECT 815.015 84.330 818.385 84.630 ;
        RECT 823.265 84.425 824.570 84.805 ;
        RECT 825.270 84.425 828.570 84.805 ;
        RECT 829.270 84.425 832.570 84.805 ;
        RECT 833.270 84.425 834.630 84.805 ;
        RECT 836.605 84.425 838.070 84.805 ;
        RECT 838.770 84.425 842.070 84.805 ;
        RECT 842.770 84.425 846.070 84.805 ;
        RECT 846.770 84.425 847.950 84.805 ;
        RECT 861.910 84.400 863.215 84.780 ;
        RECT 867.915 84.400 871.215 84.780 ;
        RECT 871.915 84.400 873.275 84.780 ;
        RECT 875.250 84.400 876.715 84.780 ;
        RECT 877.415 84.400 880.715 84.780 ;
        RECT 885.415 84.400 886.595 84.780 ;
        RECT 824.730 84.080 825.110 84.115 ;
        RECT 806.765 83.595 807.145 83.975 ;
        RECT 809.170 83.610 810.950 83.900 ;
        RECT 812.425 83.700 813.615 83.985 ;
        RECT 816.545 83.580 817.855 83.900 ;
        RECT 824.465 83.770 827.475 84.080 ;
        RECT 824.730 83.735 825.110 83.770 ;
        RECT 828.730 83.735 829.820 84.115 ;
        RECT 832.730 84.110 833.110 84.115 ;
        RECT 830.250 83.745 833.115 84.110 ;
        RECT 838.230 84.090 838.610 84.115 ;
        RECT 838.215 83.770 840.360 84.090 ;
        RECT 832.730 83.735 833.110 83.745 ;
        RECT 838.230 83.735 838.610 83.770 ;
        RECT 841.275 83.735 842.610 84.115 ;
        RECT 846.230 84.095 846.610 84.115 ;
        RECT 843.765 83.775 846.675 84.095 ;
        RECT 863.375 84.055 863.755 84.090 ;
        RECT 846.230 83.735 846.610 83.775 ;
        RECT 863.110 83.745 866.120 84.055 ;
        RECT 863.375 83.710 863.755 83.745 ;
        RECT 867.375 83.710 868.465 84.090 ;
        RECT 871.375 84.085 871.755 84.090 ;
        RECT 868.895 83.720 871.760 84.085 ;
        RECT 876.875 84.065 877.255 84.090 ;
        RECT 876.860 83.745 879.005 84.065 ;
        RECT 871.375 83.710 871.755 83.720 ;
        RECT 876.875 83.710 877.255 83.745 ;
        RECT 879.920 83.710 881.255 84.090 ;
        RECT 884.875 84.070 885.255 84.090 ;
        RECT 882.410 83.750 885.320 84.070 ;
        RECT 884.875 83.710 885.255 83.750 ;
        RECT 889.505 83.570 889.885 83.950 ;
        RECT 891.910 83.585 893.690 83.875 ;
        RECT 895.165 83.675 896.355 83.960 ;
        RECT 899.285 83.555 900.595 83.875 ;
        RECT 807.900 82.995 808.280 83.375 ;
        RECT 811.645 83.035 812.025 83.415 ;
        RECT 814.355 83.025 814.735 83.405 ;
        RECT 815.765 82.870 818.945 83.190 ;
        RECT 890.640 82.970 891.020 83.350 ;
        RECT 894.385 83.010 894.765 83.390 ;
        RECT 897.095 83.000 897.475 83.380 ;
        RECT 898.505 82.845 901.685 83.165 ;
        RECT 823.080 82.425 824.570 82.805 ;
        RECT 825.270 82.425 826.555 82.805 ;
        RECT 844.585 82.425 846.070 82.805 ;
        RECT 846.770 82.425 847.845 82.805 ;
        RECT 861.725 82.400 863.215 82.780 ;
        RECT 885.415 82.400 886.490 82.780 ;
        RECT 824.730 81.735 825.820 82.115 ;
        RECT 826.775 81.745 828.295 82.105 ;
        RECT 829.215 81.740 842.065 82.075 ;
        RECT 846.230 82.070 846.610 82.115 ;
        RECT 845.495 81.770 846.805 82.070 ;
        RECT 846.230 81.735 846.610 81.770 ;
        RECT 863.375 81.710 864.465 82.090 ;
        RECT 865.420 81.720 866.940 82.080 ;
        RECT 867.860 81.715 880.710 82.050 ;
        RECT 884.875 82.045 885.255 82.090 ;
        RECT 884.140 81.745 885.450 82.045 ;
        RECT 884.875 81.710 885.255 81.745 ;
        RECT 821.585 81.215 854.665 81.225 ;
        RECT 821.585 80.875 886.885 81.215 ;
        RECT 853.935 80.850 886.885 80.875 ;
        RECT 888.680 80.840 892.940 81.195 ;
        RECT 805.695 80.280 809.790 80.285 ;
        RECT 789.115 80.275 794.330 80.280 ;
        RECT 804.575 80.275 809.790 80.280 ;
        RECT 820.035 80.275 860.285 80.280 ;
        RECT 707.555 80.255 711.650 80.260 ;
        RECT 592.775 80.250 696.190 80.255 ;
        RECT 706.435 80.250 711.650 80.255 ;
        RECT 592.775 79.380 721.465 80.250 ;
        RECT 663.890 79.355 721.465 79.380 ;
        RECT 752.815 79.375 779.470 80.275 ;
        RECT 789.115 80.255 860.285 80.275 ;
        RECT 886.885 80.255 892.530 80.260 ;
        RECT 903.145 80.255 903.525 86.085 ;
        RECT 912.025 86.035 916.525 86.345 ;
        RECT 988.200 86.110 992.330 86.410 ;
        RECT 907.985 85.485 914.375 85.775 ;
        RECT 907.400 84.905 923.420 85.240 ;
        RECT 972.290 85.045 978.205 85.380 ;
        RECT 975.560 85.025 978.205 85.045 ;
        RECT 906.750 84.320 909.670 84.620 ;
        RECT 913.215 84.305 916.585 84.605 ;
        RECT 952.885 84.405 956.185 84.785 ;
        RECT 956.885 84.405 960.185 84.785 ;
        RECT 966.385 84.405 969.685 84.785 ;
        RECT 970.385 84.405 973.685 84.785 ;
        RECT 904.965 83.570 905.345 83.950 ;
        RECT 907.370 83.585 909.150 83.875 ;
        RECT 910.625 83.675 911.815 83.960 ;
        RECT 914.745 83.555 916.055 83.875 ;
        RECT 906.100 82.970 906.480 83.350 ;
        RECT 909.845 83.010 910.225 83.390 ;
        RECT 912.555 83.000 912.935 83.380 ;
        RECT 913.965 82.845 917.145 83.165 ;
        RECT 952.885 82.405 954.170 82.785 ;
        RECT 972.200 82.405 973.685 82.785 ;
        RECT 904.245 81.760 908.395 82.030 ;
        RECT 954.390 81.725 955.910 82.085 ;
        RECT 985.825 80.280 986.205 86.110 ;
        RECT 994.705 86.060 999.205 86.370 ;
        RECT 1003.660 86.110 1007.790 86.410 ;
        RECT 990.665 85.510 997.055 85.800 ;
        RECT 990.080 84.930 1000.735 85.265 ;
        RECT 989.430 84.345 992.350 84.645 ;
        RECT 995.895 84.330 999.265 84.630 ;
        RECT 987.645 83.595 988.025 83.975 ;
        RECT 990.050 83.610 991.830 83.900 ;
        RECT 993.305 83.700 994.495 83.985 ;
        RECT 997.425 83.580 998.735 83.900 ;
        RECT 988.780 82.995 989.160 83.375 ;
        RECT 992.525 83.035 992.905 83.415 ;
        RECT 995.235 83.025 995.615 83.405 ;
        RECT 996.645 82.870 999.825 83.190 ;
        RECT 986.575 80.280 990.670 80.285 ;
        RECT 1001.285 80.280 1001.665 86.110 ;
        RECT 1010.165 86.060 1014.665 86.370 ;
        RECT 1101.860 86.085 1105.990 86.385 ;
        RECT 1017.395 85.875 1053.305 85.900 ;
        RECT 1006.125 85.510 1012.515 85.800 ;
        RECT 1017.395 85.630 1084.645 85.875 ;
        RECT 1052.900 85.605 1084.645 85.630 ;
        RECT 1088.865 85.485 1095.255 85.775 ;
        RECT 1005.540 84.930 1016.045 85.265 ;
        RECT 1041.015 85.065 1051.565 85.400 ;
        RECT 1088.280 84.905 1098.760 85.240 ;
        RECT 1004.890 84.345 1007.810 84.645 ;
        RECT 1011.355 84.330 1014.725 84.630 ;
        RECT 1019.605 84.425 1020.910 84.805 ;
        RECT 1021.610 84.425 1024.910 84.805 ;
        RECT 1025.610 84.425 1028.910 84.805 ;
        RECT 1029.610 84.425 1030.970 84.805 ;
        RECT 1032.945 84.425 1034.410 84.805 ;
        RECT 1035.110 84.425 1038.410 84.805 ;
        RECT 1039.110 84.425 1042.410 84.805 ;
        RECT 1043.110 84.425 1044.290 84.805 ;
        RECT 1058.250 84.400 1059.555 84.780 ;
        RECT 1064.255 84.400 1067.555 84.780 ;
        RECT 1068.255 84.400 1069.615 84.780 ;
        RECT 1071.590 84.400 1073.055 84.780 ;
        RECT 1073.755 84.400 1077.055 84.780 ;
        RECT 1081.755 84.400 1082.935 84.780 ;
        RECT 1021.070 84.080 1021.450 84.115 ;
        RECT 1003.105 83.595 1003.485 83.975 ;
        RECT 1005.510 83.610 1007.290 83.900 ;
        RECT 1008.765 83.700 1009.955 83.985 ;
        RECT 1012.885 83.580 1014.195 83.900 ;
        RECT 1020.805 83.770 1023.815 84.080 ;
        RECT 1021.070 83.735 1021.450 83.770 ;
        RECT 1025.070 83.735 1026.160 84.115 ;
        RECT 1029.070 84.110 1029.450 84.115 ;
        RECT 1026.590 83.745 1029.455 84.110 ;
        RECT 1034.570 84.090 1034.950 84.115 ;
        RECT 1034.555 83.770 1036.700 84.090 ;
        RECT 1029.070 83.735 1029.450 83.745 ;
        RECT 1034.570 83.735 1034.950 83.770 ;
        RECT 1037.615 83.735 1038.950 84.115 ;
        RECT 1042.570 84.095 1042.950 84.115 ;
        RECT 1040.105 83.775 1043.015 84.095 ;
        RECT 1059.715 84.055 1060.095 84.090 ;
        RECT 1042.570 83.735 1042.950 83.775 ;
        RECT 1059.450 83.745 1062.460 84.055 ;
        RECT 1059.715 83.710 1060.095 83.745 ;
        RECT 1063.715 83.710 1064.805 84.090 ;
        RECT 1067.715 84.085 1068.095 84.090 ;
        RECT 1065.235 83.720 1068.100 84.085 ;
        RECT 1073.215 84.065 1073.595 84.090 ;
        RECT 1073.200 83.745 1075.345 84.065 ;
        RECT 1067.715 83.710 1068.095 83.720 ;
        RECT 1073.215 83.710 1073.595 83.745 ;
        RECT 1076.260 83.710 1077.595 84.090 ;
        RECT 1081.215 84.070 1081.595 84.090 ;
        RECT 1078.750 83.750 1081.660 84.070 ;
        RECT 1081.215 83.710 1081.595 83.750 ;
        RECT 1085.845 83.570 1086.225 83.950 ;
        RECT 1088.250 83.585 1090.030 83.875 ;
        RECT 1091.505 83.675 1092.695 83.960 ;
        RECT 1095.625 83.555 1096.935 83.875 ;
        RECT 1004.240 82.995 1004.620 83.375 ;
        RECT 1007.985 83.035 1008.365 83.415 ;
        RECT 1010.695 83.025 1011.075 83.405 ;
        RECT 1012.105 82.870 1015.285 83.190 ;
        RECT 1086.980 82.970 1087.360 83.350 ;
        RECT 1090.725 83.010 1091.105 83.390 ;
        RECT 1093.435 83.000 1093.815 83.380 ;
        RECT 1094.845 82.845 1098.025 83.165 ;
        RECT 1019.420 82.425 1020.910 82.805 ;
        RECT 1021.610 82.425 1022.895 82.805 ;
        RECT 1040.925 82.425 1042.410 82.805 ;
        RECT 1043.110 82.425 1044.185 82.805 ;
        RECT 1058.065 82.400 1059.555 82.780 ;
        RECT 1081.755 82.400 1082.830 82.780 ;
        RECT 1021.070 81.735 1022.160 82.115 ;
        RECT 1023.115 81.745 1024.635 82.105 ;
        RECT 1025.555 81.740 1038.405 82.075 ;
        RECT 1042.570 82.070 1042.950 82.115 ;
        RECT 1041.835 81.770 1043.145 82.070 ;
        RECT 1042.570 81.735 1042.950 81.770 ;
        RECT 1059.715 81.710 1060.805 82.090 ;
        RECT 1061.760 81.720 1063.280 82.080 ;
        RECT 1064.200 81.715 1077.050 82.050 ;
        RECT 1081.215 82.045 1081.595 82.090 ;
        RECT 1080.480 81.745 1081.790 82.045 ;
        RECT 1081.215 81.710 1081.595 81.745 ;
        RECT 1017.925 81.215 1051.005 81.225 ;
        RECT 1017.925 80.875 1083.225 81.215 ;
        RECT 1050.275 80.850 1083.225 80.875 ;
        RECT 1085.020 80.840 1089.280 81.195 ;
        RECT 1002.035 80.280 1006.130 80.285 ;
        RECT 985.455 80.275 990.670 80.280 ;
        RECT 1000.915 80.275 1006.130 80.280 ;
        RECT 1016.375 80.275 1056.625 80.280 ;
        RECT 903.895 80.255 907.990 80.260 ;
        RECT 789.115 80.250 892.530 80.255 ;
        RECT 902.775 80.250 907.990 80.255 ;
        RECT 789.115 79.380 917.805 80.250 ;
        RECT 860.230 79.355 917.805 79.380 ;
        RECT 949.200 79.360 975.855 80.260 ;
        RECT 985.455 80.255 1056.625 80.275 ;
        RECT 1083.225 80.255 1088.870 80.260 ;
        RECT 1099.485 80.255 1099.865 86.085 ;
        RECT 1108.365 86.035 1112.865 86.345 ;
        RECT 1184.540 86.110 1188.670 86.410 ;
        RECT 1104.325 85.485 1110.715 85.775 ;
        RECT 1103.740 84.905 1119.760 85.240 ;
        RECT 1168.615 85.050 1174.530 85.385 ;
        RECT 1171.885 85.030 1174.530 85.050 ;
        RECT 1103.090 84.320 1106.010 84.620 ;
        RECT 1109.555 84.305 1112.925 84.605 ;
        RECT 1149.210 84.410 1152.510 84.790 ;
        RECT 1153.210 84.410 1156.510 84.790 ;
        RECT 1162.710 84.410 1166.010 84.790 ;
        RECT 1166.710 84.410 1170.010 84.790 ;
        RECT 1101.305 83.570 1101.685 83.950 ;
        RECT 1103.710 83.585 1105.490 83.875 ;
        RECT 1106.965 83.675 1108.155 83.960 ;
        RECT 1111.085 83.555 1112.395 83.875 ;
        RECT 1102.440 82.970 1102.820 83.350 ;
        RECT 1106.185 83.010 1106.565 83.390 ;
        RECT 1108.895 83.000 1109.275 83.380 ;
        RECT 1110.305 82.845 1113.485 83.165 ;
        RECT 1149.210 82.410 1150.495 82.790 ;
        RECT 1168.525 82.410 1170.010 82.790 ;
        RECT 1100.585 81.760 1104.735 82.030 ;
        RECT 1150.715 81.730 1152.235 82.090 ;
        RECT 1182.165 80.280 1182.545 86.110 ;
        RECT 1191.045 86.060 1195.545 86.370 ;
        RECT 1200.000 86.110 1204.130 86.410 ;
        RECT 1187.005 85.510 1193.395 85.800 ;
        RECT 1186.420 84.930 1197.075 85.265 ;
        RECT 1185.770 84.345 1188.690 84.645 ;
        RECT 1192.235 84.330 1195.605 84.630 ;
        RECT 1183.985 83.595 1184.365 83.975 ;
        RECT 1186.390 83.610 1188.170 83.900 ;
        RECT 1189.645 83.700 1190.835 83.985 ;
        RECT 1193.765 83.580 1195.075 83.900 ;
        RECT 1185.120 82.995 1185.500 83.375 ;
        RECT 1188.865 83.035 1189.245 83.415 ;
        RECT 1191.575 83.025 1191.955 83.405 ;
        RECT 1192.985 82.870 1196.165 83.190 ;
        RECT 1182.915 80.280 1187.010 80.285 ;
        RECT 1197.625 80.280 1198.005 86.110 ;
        RECT 1206.505 86.060 1211.005 86.370 ;
        RECT 1282.740 86.085 1286.870 86.385 ;
        RECT 1289.245 86.035 1293.745 86.345 ;
        RECT 1298.200 86.085 1302.330 86.385 ;
        RECT 1213.735 85.875 1249.645 85.900 ;
        RECT 1202.465 85.510 1208.855 85.800 ;
        RECT 1213.735 85.630 1280.985 85.875 ;
        RECT 1249.240 85.605 1280.985 85.630 ;
        RECT 1285.205 85.485 1291.595 85.775 ;
        RECT 1201.880 84.930 1212.385 85.265 ;
        RECT 1237.355 85.065 1247.905 85.400 ;
        RECT 1276.000 85.040 1279.945 85.375 ;
        RECT 1284.620 84.905 1295.100 85.240 ;
        RECT 1201.230 84.345 1204.150 84.645 ;
        RECT 1207.695 84.330 1211.065 84.630 ;
        RECT 1215.945 84.425 1217.250 84.805 ;
        RECT 1217.950 84.425 1221.250 84.805 ;
        RECT 1221.950 84.425 1225.250 84.805 ;
        RECT 1225.950 84.425 1227.310 84.805 ;
        RECT 1229.285 84.425 1230.750 84.805 ;
        RECT 1231.450 84.425 1234.750 84.805 ;
        RECT 1235.450 84.425 1238.750 84.805 ;
        RECT 1239.450 84.425 1240.630 84.805 ;
        RECT 1254.590 84.400 1255.895 84.780 ;
        RECT 1256.595 84.400 1259.895 84.780 ;
        RECT 1260.595 84.400 1263.895 84.780 ;
        RECT 1264.595 84.400 1265.955 84.780 ;
        RECT 1267.930 84.400 1269.395 84.780 ;
        RECT 1270.095 84.400 1273.395 84.780 ;
        RECT 1274.095 84.400 1277.395 84.780 ;
        RECT 1278.095 84.400 1279.275 84.780 ;
        RECT 1283.970 84.320 1286.890 84.620 ;
        RECT 1290.435 84.305 1293.805 84.605 ;
        RECT 1217.410 84.080 1217.790 84.115 ;
        RECT 1199.445 83.595 1199.825 83.975 ;
        RECT 1201.850 83.610 1203.630 83.900 ;
        RECT 1205.105 83.700 1206.295 83.985 ;
        RECT 1209.225 83.580 1210.535 83.900 ;
        RECT 1217.145 83.770 1220.155 84.080 ;
        RECT 1217.410 83.735 1217.790 83.770 ;
        RECT 1221.410 83.735 1222.500 84.115 ;
        RECT 1225.410 84.110 1225.790 84.115 ;
        RECT 1222.930 83.745 1225.795 84.110 ;
        RECT 1230.910 84.090 1231.290 84.115 ;
        RECT 1230.895 83.770 1233.040 84.090 ;
        RECT 1225.410 83.735 1225.790 83.745 ;
        RECT 1230.910 83.735 1231.290 83.770 ;
        RECT 1233.955 83.735 1235.290 84.115 ;
        RECT 1238.910 84.095 1239.290 84.115 ;
        RECT 1236.445 83.775 1239.355 84.095 ;
        RECT 1256.055 84.055 1256.435 84.090 ;
        RECT 1238.910 83.735 1239.290 83.775 ;
        RECT 1255.790 83.745 1258.800 84.055 ;
        RECT 1256.055 83.710 1256.435 83.745 ;
        RECT 1260.055 83.710 1261.145 84.090 ;
        RECT 1264.055 84.085 1264.435 84.090 ;
        RECT 1261.575 83.720 1264.440 84.085 ;
        RECT 1269.555 84.065 1269.935 84.090 ;
        RECT 1269.540 83.745 1271.685 84.065 ;
        RECT 1264.055 83.710 1264.435 83.720 ;
        RECT 1269.555 83.710 1269.935 83.745 ;
        RECT 1272.600 83.710 1273.935 84.090 ;
        RECT 1277.555 84.070 1277.935 84.090 ;
        RECT 1275.090 83.750 1278.000 84.070 ;
        RECT 1277.555 83.710 1277.935 83.750 ;
        RECT 1282.185 83.570 1282.565 83.950 ;
        RECT 1284.590 83.585 1286.370 83.875 ;
        RECT 1287.845 83.675 1289.035 83.960 ;
        RECT 1291.965 83.555 1293.275 83.875 ;
        RECT 1200.580 82.995 1200.960 83.375 ;
        RECT 1204.325 83.035 1204.705 83.415 ;
        RECT 1207.035 83.025 1207.415 83.405 ;
        RECT 1208.445 82.870 1211.625 83.190 ;
        RECT 1283.320 82.970 1283.700 83.350 ;
        RECT 1287.065 83.010 1287.445 83.390 ;
        RECT 1289.775 83.000 1290.155 83.380 ;
        RECT 1291.185 82.845 1294.365 83.165 ;
        RECT 1215.760 82.425 1217.250 82.805 ;
        RECT 1217.950 82.425 1219.235 82.805 ;
        RECT 1237.265 82.425 1238.750 82.805 ;
        RECT 1239.450 82.425 1240.525 82.805 ;
        RECT 1254.405 82.400 1255.895 82.780 ;
        RECT 1256.595 82.400 1257.880 82.780 ;
        RECT 1275.910 82.400 1277.395 82.780 ;
        RECT 1278.095 82.400 1279.170 82.780 ;
        RECT 1217.410 81.735 1218.500 82.115 ;
        RECT 1219.455 81.745 1220.975 82.105 ;
        RECT 1221.895 81.740 1234.745 82.075 ;
        RECT 1238.910 82.070 1239.290 82.115 ;
        RECT 1238.175 81.770 1239.485 82.070 ;
        RECT 1238.910 81.735 1239.290 81.770 ;
        RECT 1256.055 81.710 1257.145 82.090 ;
        RECT 1258.100 81.720 1259.620 82.080 ;
        RECT 1260.540 81.715 1273.390 82.050 ;
        RECT 1277.555 82.045 1277.935 82.090 ;
        RECT 1276.820 81.745 1278.130 82.045 ;
        RECT 1277.555 81.710 1277.935 81.745 ;
        RECT 1214.265 81.215 1247.345 81.225 ;
        RECT 1214.265 80.875 1279.565 81.215 ;
        RECT 1246.615 80.850 1279.565 80.875 ;
        RECT 1281.360 80.840 1285.620 81.195 ;
        RECT 1198.375 80.280 1202.470 80.285 ;
        RECT 1181.795 80.275 1187.010 80.280 ;
        RECT 1197.255 80.275 1202.470 80.280 ;
        RECT 1212.715 80.275 1252.965 80.280 ;
        RECT 1100.235 80.255 1104.330 80.260 ;
        RECT 985.455 80.250 1088.870 80.255 ;
        RECT 1099.115 80.250 1104.330 80.255 ;
        RECT 985.455 79.380 1114.145 80.250 ;
        RECT 1056.570 79.355 1114.145 79.380 ;
        RECT 1145.525 79.365 1172.180 80.265 ;
        RECT 1181.795 80.255 1252.965 80.275 ;
        RECT 1279.565 80.255 1285.210 80.260 ;
        RECT 1295.825 80.255 1296.205 86.085 ;
        RECT 1304.705 86.035 1309.205 86.345 ;
        RECT 1300.665 85.485 1307.055 85.775 ;
        RECT 1299.430 84.320 1302.350 84.620 ;
        RECT 1305.895 84.305 1309.265 84.605 ;
        RECT 1297.645 83.570 1298.025 83.950 ;
        RECT 1303.305 83.675 1304.495 83.960 ;
        RECT 1302.525 83.010 1302.905 83.390 ;
        RECT 1306.645 82.845 1309.825 83.165 ;
        RECT 1296.925 81.760 1301.075 82.030 ;
        RECT 1296.575 80.255 1300.670 80.260 ;
        RECT 1181.795 80.250 1285.210 80.255 ;
        RECT 1295.455 80.250 1300.670 80.255 ;
        RECT 1181.795 79.380 1310.485 80.250 ;
        RECT 1252.910 79.355 1310.485 79.380 ;
        RECT 467.515 79.320 525.090 79.345 ;
        RECT 76.075 75.560 132.430 75.580 ;
        RECT 272.440 75.560 328.795 75.580 ;
        RECT -81.605 74.470 -56.170 75.370 ;
        RECT -31.280 74.550 -5.845 75.450 ;
        RECT 3.765 74.680 132.430 75.560 ;
        RECT 3.765 74.660 76.155 74.680 ;
        RECT -79.120 72.290 -77.920 72.670 ;
        RECT -76.165 72.075 -73.890 72.585 ;
        RECT -71.265 72.075 -68.965 72.585 ;
        RECT -66.670 72.075 -64.390 72.585 ;
        RECT -59.595 72.390 -58.360 72.770 ;
        RECT -28.795 72.370 -27.595 72.750 ;
        RECT -25.840 72.155 -23.565 72.665 ;
        RECT -20.940 72.155 -18.640 72.665 ;
        RECT -16.345 72.155 -14.065 72.665 ;
        RECT -9.270 72.470 -8.035 72.850 ;
        RECT -79.120 69.990 -75.860 70.370 ;
        RECT -75.120 69.990 -71.860 70.370 ;
        RECT -65.620 69.990 -62.360 70.370 ;
        RECT -61.620 69.990 -58.360 70.370 ;
        RECT -28.795 70.070 -25.535 70.450 ;
        RECT -24.795 70.070 -21.535 70.450 ;
        RECT -15.295 70.070 -12.035 70.450 ;
        RECT -11.295 70.070 -8.035 70.450 ;
        RECT -78.455 68.405 -56.170 68.415 ;
        RECT -78.455 68.075 -54.630 68.405 ;
        RECT -28.130 68.155 -1.835 68.495 ;
        RECT -56.390 68.055 -54.630 68.075 ;
        RECT 4.135 67.500 4.515 74.660 ;
        RECT 5.965 70.445 9.340 70.845 ;
        RECT 9.710 70.205 10.090 70.585 ;
        RECT 12.425 70.245 12.805 70.625 ;
        RECT 16.610 70.195 16.990 70.575 ;
        RECT 7.035 69.780 8.775 70.070 ;
        RECT 10.825 69.730 12.025 70.020 ;
        RECT 13.535 69.700 16.145 70.125 ;
        RECT 17.745 69.795 18.125 70.175 ;
        RECT 5.280 69.020 18.845 69.335 ;
        RECT 5.275 68.275 18.835 68.575 ;
        RECT 5.295 67.560 12.020 67.860 ;
        RECT 15.720 67.260 18.825 67.535 ;
        RECT 19.595 67.500 19.975 74.660 ;
        RECT 73.060 73.675 101.835 73.695 ;
        RECT 36.235 73.410 101.835 73.675 ;
        RECT 36.235 73.390 73.785 73.410 ;
        RECT 103.505 73.390 110.210 73.690 ;
        RECT 37.745 72.480 39.200 72.860 ;
        RECT 39.940 72.480 41.140 72.860 ;
        RECT 42.895 72.265 45.170 72.775 ;
        RECT 47.795 72.265 50.095 72.775 ;
        RECT 52.390 72.265 54.670 72.775 ;
        RECT 59.465 72.580 60.700 72.960 ;
        RECT 61.440 72.580 62.720 72.960 ;
        RECT 76.365 72.500 77.820 72.880 ;
        RECT 81.515 72.285 83.790 72.795 ;
        RECT 86.415 72.285 88.715 72.795 ;
        RECT 91.010 72.285 93.290 72.795 ;
        RECT 100.060 72.600 101.340 72.980 ;
        RECT 60.880 72.225 61.260 72.260 ;
        RECT 99.500 72.245 99.880 72.280 ;
        RECT 39.380 72.120 39.760 72.160 ;
        RECT 39.310 71.815 42.145 72.120 ;
        RECT 58.125 71.915 61.260 72.225 ;
        RECT 78.000 72.140 78.380 72.180 ;
        RECT 60.880 71.880 61.260 71.915 ;
        RECT 77.930 71.835 80.765 72.140 ;
        RECT 96.745 71.935 99.880 72.245 ;
        RECT 99.500 71.900 99.880 71.935 ;
        RECT 39.380 71.780 39.760 71.815 ;
        RECT 78.000 71.800 78.380 71.835 ;
        RECT 21.425 70.405 24.830 70.845 ;
        RECT 25.170 70.205 25.550 70.585 ;
        RECT 27.885 70.245 28.265 70.625 ;
        RECT 32.070 70.195 32.450 70.575 ;
        RECT 37.905 70.180 39.200 70.560 ;
        RECT 39.940 70.180 43.200 70.560 ;
        RECT 43.940 70.180 47.200 70.560 ;
        RECT 47.940 70.180 49.125 70.560 ;
        RECT 51.390 70.180 52.700 70.560 ;
        RECT 53.440 70.180 56.700 70.560 ;
        RECT 57.440 70.180 60.700 70.560 ;
        RECT 61.440 70.180 62.455 70.560 ;
        RECT 76.525 70.200 77.820 70.580 ;
        RECT 82.560 70.200 85.820 70.580 ;
        RECT 86.560 70.200 87.745 70.580 ;
        RECT 90.010 70.200 91.320 70.580 ;
        RECT 92.060 70.200 95.320 70.580 ;
        RECT 100.060 70.200 101.075 70.580 ;
        RECT 104.140 70.445 107.555 70.865 ;
        RECT 107.885 70.225 108.265 70.605 ;
        RECT 110.600 70.265 110.980 70.645 ;
        RECT 114.785 70.215 115.165 70.595 ;
        RECT 22.495 69.780 24.235 70.070 ;
        RECT 26.285 69.730 27.485 70.020 ;
        RECT 28.995 69.700 31.590 70.075 ;
        RECT 33.205 69.795 33.585 70.175 ;
        RECT 39.380 69.480 39.760 69.860 ;
        RECT 43.380 69.480 43.760 69.860 ;
        RECT 47.380 69.815 47.760 69.860 ;
        RECT 52.880 69.815 53.260 69.860 ;
        RECT 47.330 69.500 53.265 69.815 ;
        RECT 47.380 69.480 47.760 69.500 ;
        RECT 52.880 69.480 53.260 69.500 ;
        RECT 56.880 69.480 57.260 69.860 ;
        RECT 60.880 69.480 61.260 69.860 ;
        RECT 78.000 69.500 78.380 69.880 ;
        RECT 82.000 69.500 82.380 69.880 ;
        RECT 86.000 69.835 86.380 69.880 ;
        RECT 91.500 69.835 91.880 69.880 ;
        RECT 85.950 69.520 91.885 69.835 ;
        RECT 86.000 69.500 86.380 69.520 ;
        RECT 91.500 69.500 91.880 69.520 ;
        RECT 95.500 69.500 95.880 69.880 ;
        RECT 99.500 69.500 99.880 69.880 ;
        RECT 105.210 69.800 106.950 70.090 ;
        RECT 109.000 69.750 110.200 70.040 ;
        RECT 111.710 69.710 114.340 70.165 ;
        RECT 115.920 69.815 116.300 70.195 ;
        RECT 20.735 69.020 34.560 69.320 ;
        RECT 36.235 68.855 52.245 69.230 ;
        RECT 70.090 68.875 90.865 69.250 ;
        RECT 20.740 68.275 39.160 68.575 ;
        RECT 40.605 68.265 67.915 68.605 ;
        RECT 20.220 67.560 27.480 67.860 ;
        RECT 5.275 66.940 9.400 67.210 ;
        RECT 20.775 67.025 24.860 67.295 ;
        RECT 31.180 67.260 34.930 67.535 ;
        RECT 36.235 67.500 62.465 67.890 ;
        RECT 69.120 67.520 101.085 67.910 ;
        RECT 113.895 67.280 117.025 67.555 ;
        RECT 117.770 67.520 118.150 74.680 ;
        RECT 164.890 74.560 190.325 75.460 ;
        RECT 200.130 74.680 328.795 75.560 ;
        RECT 665.215 75.545 721.570 75.565 ;
        RECT 861.555 75.545 917.910 75.565 ;
        RECT 1057.895 75.545 1114.250 75.565 ;
        RECT 1254.235 75.545 1310.590 75.565 ;
        RECT 468.840 75.510 525.195 75.530 ;
        RECT 200.130 74.660 272.520 74.680 ;
        RECT 119.010 72.220 125.750 72.520 ;
        RECT 167.375 72.380 168.575 72.760 ;
        RECT 170.330 72.165 172.605 72.675 ;
        RECT 175.230 72.165 177.530 72.675 ;
        RECT 179.825 72.165 182.105 72.675 ;
        RECT 186.900 72.480 188.135 72.860 ;
        RECT 119.600 70.425 123.055 70.865 ;
        RECT 123.345 70.225 123.725 70.605 ;
        RECT 126.060 70.265 126.440 70.645 ;
        RECT 130.245 70.215 130.625 70.595 ;
        RECT 120.670 69.800 122.410 70.090 ;
        RECT 124.460 69.750 125.660 70.040 ;
        RECT 127.170 69.720 129.795 70.130 ;
        RECT 131.380 69.815 131.760 70.195 ;
        RECT 167.375 70.080 170.635 70.460 ;
        RECT 171.375 70.080 174.635 70.460 ;
        RECT 180.875 70.080 184.135 70.460 ;
        RECT 184.875 70.080 188.135 70.460 ;
        RECT 118.415 69.040 134.335 69.340 ;
        RECT 118.950 68.295 135.895 68.595 ;
        RECT 168.040 68.165 194.335 68.505 ;
        RECT 129.355 67.280 137.055 67.555 ;
        RECT 200.500 67.500 200.880 74.660 ;
        RECT 202.330 70.445 205.705 70.845 ;
        RECT 206.075 70.205 206.455 70.585 ;
        RECT 208.790 70.245 209.170 70.625 ;
        RECT 212.975 70.195 213.355 70.575 ;
        RECT 203.400 69.780 205.140 70.070 ;
        RECT 207.190 69.730 208.390 70.020 ;
        RECT 209.900 69.700 212.510 70.125 ;
        RECT 214.110 69.795 214.490 70.175 ;
        RECT 201.645 69.020 215.210 69.335 ;
        RECT 201.640 68.275 215.200 68.575 ;
        RECT 201.660 67.560 208.385 67.860 ;
        RECT 212.085 67.260 215.190 67.535 ;
        RECT 215.960 67.500 216.340 74.660 ;
        RECT 269.425 73.675 298.200 73.695 ;
        RECT 232.600 73.410 298.200 73.675 ;
        RECT 232.600 73.390 270.150 73.410 ;
        RECT 299.870 73.390 306.575 73.690 ;
        RECT 234.110 72.480 235.565 72.860 ;
        RECT 236.305 72.480 237.505 72.860 ;
        RECT 239.260 72.265 241.535 72.775 ;
        RECT 244.160 72.265 246.460 72.775 ;
        RECT 248.755 72.265 251.035 72.775 ;
        RECT 255.830 72.580 257.065 72.960 ;
        RECT 257.805 72.580 259.085 72.960 ;
        RECT 272.730 72.500 274.185 72.880 ;
        RECT 277.880 72.285 280.155 72.795 ;
        RECT 282.780 72.285 285.080 72.795 ;
        RECT 287.375 72.285 289.655 72.795 ;
        RECT 296.425 72.600 297.705 72.980 ;
        RECT 257.245 72.225 257.625 72.260 ;
        RECT 295.865 72.245 296.245 72.280 ;
        RECT 235.745 72.120 236.125 72.160 ;
        RECT 235.675 71.815 238.510 72.120 ;
        RECT 254.490 71.915 257.625 72.225 ;
        RECT 274.365 72.140 274.745 72.180 ;
        RECT 257.245 71.880 257.625 71.915 ;
        RECT 274.295 71.835 277.130 72.140 ;
        RECT 293.110 71.935 296.245 72.245 ;
        RECT 295.865 71.900 296.245 71.935 ;
        RECT 235.745 71.780 236.125 71.815 ;
        RECT 274.365 71.800 274.745 71.835 ;
        RECT 217.790 70.405 221.195 70.845 ;
        RECT 221.535 70.205 221.915 70.585 ;
        RECT 224.250 70.245 224.630 70.625 ;
        RECT 228.435 70.195 228.815 70.575 ;
        RECT 234.270 70.180 235.565 70.560 ;
        RECT 236.305 70.180 239.565 70.560 ;
        RECT 240.305 70.180 243.565 70.560 ;
        RECT 244.305 70.180 245.490 70.560 ;
        RECT 247.755 70.180 249.065 70.560 ;
        RECT 249.805 70.180 253.065 70.560 ;
        RECT 253.805 70.180 257.065 70.560 ;
        RECT 257.805 70.180 258.820 70.560 ;
        RECT 272.890 70.200 274.185 70.580 ;
        RECT 278.925 70.200 282.185 70.580 ;
        RECT 282.925 70.200 284.110 70.580 ;
        RECT 286.375 70.200 287.685 70.580 ;
        RECT 288.425 70.200 291.685 70.580 ;
        RECT 296.425 70.200 297.440 70.580 ;
        RECT 300.505 70.445 303.920 70.865 ;
        RECT 304.250 70.225 304.630 70.605 ;
        RECT 306.965 70.265 307.345 70.645 ;
        RECT 311.150 70.215 311.530 70.595 ;
        RECT 218.860 69.780 220.600 70.070 ;
        RECT 222.650 69.730 223.850 70.020 ;
        RECT 225.360 69.700 227.955 70.075 ;
        RECT 229.570 69.795 229.950 70.175 ;
        RECT 235.745 69.480 236.125 69.860 ;
        RECT 239.745 69.480 240.125 69.860 ;
        RECT 243.745 69.815 244.125 69.860 ;
        RECT 249.245 69.815 249.625 69.860 ;
        RECT 243.695 69.500 249.630 69.815 ;
        RECT 243.745 69.480 244.125 69.500 ;
        RECT 249.245 69.480 249.625 69.500 ;
        RECT 253.245 69.480 253.625 69.860 ;
        RECT 257.245 69.480 257.625 69.860 ;
        RECT 274.365 69.500 274.745 69.880 ;
        RECT 278.365 69.500 278.745 69.880 ;
        RECT 282.365 69.835 282.745 69.880 ;
        RECT 287.865 69.835 288.245 69.880 ;
        RECT 282.315 69.520 288.250 69.835 ;
        RECT 282.365 69.500 282.745 69.520 ;
        RECT 287.865 69.500 288.245 69.520 ;
        RECT 291.865 69.500 292.245 69.880 ;
        RECT 295.865 69.500 296.245 69.880 ;
        RECT 301.575 69.800 303.315 70.090 ;
        RECT 305.365 69.750 306.565 70.040 ;
        RECT 308.075 69.710 310.705 70.165 ;
        RECT 312.285 69.815 312.665 70.195 ;
        RECT 217.100 69.020 230.925 69.320 ;
        RECT 232.600 68.855 248.610 69.230 ;
        RECT 266.455 68.875 287.230 69.250 ;
        RECT 217.105 68.275 235.525 68.575 ;
        RECT 236.970 68.265 264.280 68.605 ;
        RECT 216.585 67.560 223.845 67.860 ;
        RECT 65.965 67.155 93.525 67.165 ;
        RECT 36.235 67.135 54.905 67.145 ;
        RECT 65.965 67.135 102.530 67.155 ;
        RECT 36.235 66.845 102.530 67.135 ;
        RECT 201.640 66.940 205.765 67.210 ;
        RECT 217.140 67.025 221.225 67.295 ;
        RECT 227.545 67.260 231.295 67.535 ;
        RECT 232.600 67.500 258.830 67.890 ;
        RECT 265.485 67.520 297.450 67.910 ;
        RECT 310.260 67.280 313.390 67.555 ;
        RECT 314.135 67.520 314.515 74.680 ;
        RECT 361.280 74.520 386.715 75.420 ;
        RECT 396.530 74.630 525.195 75.510 ;
        RECT 396.530 74.610 468.920 74.630 ;
        RECT 315.375 72.220 322.115 72.520 ;
        RECT 363.765 72.340 364.965 72.720 ;
        RECT 366.720 72.125 368.995 72.635 ;
        RECT 371.620 72.125 373.920 72.635 ;
        RECT 376.215 72.125 378.495 72.635 ;
        RECT 383.290 72.440 384.525 72.820 ;
        RECT 315.965 70.425 319.420 70.865 ;
        RECT 319.710 70.225 320.090 70.605 ;
        RECT 322.425 70.265 322.805 70.645 ;
        RECT 326.610 70.215 326.990 70.595 ;
        RECT 317.035 69.800 318.775 70.090 ;
        RECT 320.825 69.750 322.025 70.040 ;
        RECT 323.535 69.720 326.160 70.130 ;
        RECT 327.745 69.815 328.125 70.195 ;
        RECT 363.765 70.040 367.025 70.420 ;
        RECT 367.765 70.040 371.025 70.420 ;
        RECT 377.265 70.040 380.525 70.420 ;
        RECT 381.265 70.040 384.525 70.420 ;
        RECT 314.780 69.040 330.700 69.340 ;
        RECT 315.315 68.295 332.260 68.595 ;
        RECT 364.430 68.125 390.725 68.465 ;
        RECT 325.720 67.280 333.420 67.555 ;
        RECT 396.900 67.450 397.280 74.610 ;
        RECT 398.730 70.395 402.105 70.795 ;
        RECT 402.475 70.155 402.855 70.535 ;
        RECT 405.190 70.195 405.570 70.575 ;
        RECT 409.375 70.145 409.755 70.525 ;
        RECT 399.800 69.730 401.540 70.020 ;
        RECT 403.590 69.680 404.790 69.970 ;
        RECT 406.300 69.650 408.910 70.075 ;
        RECT 410.510 69.745 410.890 70.125 ;
        RECT 398.045 68.970 411.610 69.285 ;
        RECT 398.040 68.225 411.600 68.525 ;
        RECT 398.060 67.510 404.785 67.810 ;
        RECT 408.485 67.210 411.590 67.485 ;
        RECT 412.360 67.450 412.740 74.610 ;
        RECT 465.825 73.625 494.600 73.645 ;
        RECT 429.000 73.360 494.600 73.625 ;
        RECT 429.000 73.340 466.550 73.360 ;
        RECT 496.270 73.340 502.975 73.640 ;
        RECT 430.510 72.430 431.965 72.810 ;
        RECT 432.705 72.430 433.905 72.810 ;
        RECT 435.660 72.215 437.935 72.725 ;
        RECT 440.560 72.215 442.860 72.725 ;
        RECT 445.155 72.215 447.435 72.725 ;
        RECT 452.230 72.530 453.465 72.910 ;
        RECT 454.205 72.530 455.485 72.910 ;
        RECT 469.130 72.450 470.585 72.830 ;
        RECT 474.280 72.235 476.555 72.745 ;
        RECT 479.180 72.235 481.480 72.745 ;
        RECT 483.775 72.235 486.055 72.745 ;
        RECT 492.825 72.550 494.105 72.930 ;
        RECT 453.645 72.175 454.025 72.210 ;
        RECT 492.265 72.195 492.645 72.230 ;
        RECT 432.145 72.070 432.525 72.110 ;
        RECT 432.075 71.765 434.910 72.070 ;
        RECT 450.890 71.865 454.025 72.175 ;
        RECT 470.765 72.090 471.145 72.130 ;
        RECT 453.645 71.830 454.025 71.865 ;
        RECT 470.695 71.785 473.530 72.090 ;
        RECT 489.510 71.885 492.645 72.195 ;
        RECT 492.265 71.850 492.645 71.885 ;
        RECT 432.145 71.730 432.525 71.765 ;
        RECT 470.765 71.750 471.145 71.785 ;
        RECT 414.190 70.355 417.595 70.795 ;
        RECT 417.935 70.155 418.315 70.535 ;
        RECT 420.650 70.195 421.030 70.575 ;
        RECT 424.835 70.145 425.215 70.525 ;
        RECT 430.670 70.130 431.965 70.510 ;
        RECT 432.705 70.130 435.965 70.510 ;
        RECT 436.705 70.130 439.965 70.510 ;
        RECT 440.705 70.130 441.890 70.510 ;
        RECT 444.155 70.130 445.465 70.510 ;
        RECT 446.205 70.130 449.465 70.510 ;
        RECT 450.205 70.130 453.465 70.510 ;
        RECT 454.205 70.130 455.220 70.510 ;
        RECT 469.290 70.150 470.585 70.530 ;
        RECT 475.325 70.150 478.585 70.530 ;
        RECT 479.325 70.150 480.510 70.530 ;
        RECT 482.775 70.150 484.085 70.530 ;
        RECT 484.825 70.150 488.085 70.530 ;
        RECT 492.825 70.150 493.840 70.530 ;
        RECT 496.905 70.395 500.320 70.815 ;
        RECT 500.650 70.175 501.030 70.555 ;
        RECT 503.365 70.215 503.745 70.595 ;
        RECT 507.550 70.165 507.930 70.545 ;
        RECT 415.260 69.730 417.000 70.020 ;
        RECT 419.050 69.680 420.250 69.970 ;
        RECT 421.760 69.650 424.355 70.025 ;
        RECT 425.970 69.745 426.350 70.125 ;
        RECT 432.145 69.430 432.525 69.810 ;
        RECT 436.145 69.430 436.525 69.810 ;
        RECT 440.145 69.765 440.525 69.810 ;
        RECT 445.645 69.765 446.025 69.810 ;
        RECT 440.095 69.450 446.030 69.765 ;
        RECT 440.145 69.430 440.525 69.450 ;
        RECT 445.645 69.430 446.025 69.450 ;
        RECT 449.645 69.430 450.025 69.810 ;
        RECT 453.645 69.430 454.025 69.810 ;
        RECT 470.765 69.450 471.145 69.830 ;
        RECT 474.765 69.450 475.145 69.830 ;
        RECT 478.765 69.785 479.145 69.830 ;
        RECT 484.265 69.785 484.645 69.830 ;
        RECT 478.715 69.470 484.650 69.785 ;
        RECT 478.765 69.450 479.145 69.470 ;
        RECT 484.265 69.450 484.645 69.470 ;
        RECT 488.265 69.450 488.645 69.830 ;
        RECT 492.265 69.450 492.645 69.830 ;
        RECT 497.975 69.750 499.715 70.040 ;
        RECT 501.765 69.700 502.965 69.990 ;
        RECT 504.475 69.660 507.105 70.115 ;
        RECT 508.685 69.765 509.065 70.145 ;
        RECT 413.500 68.970 427.325 69.270 ;
        RECT 429.000 68.805 445.010 69.180 ;
        RECT 462.855 68.825 483.630 69.200 ;
        RECT 413.505 68.225 431.925 68.525 ;
        RECT 433.370 68.215 460.680 68.555 ;
        RECT 412.985 67.510 420.245 67.810 ;
        RECT 262.330 67.155 289.890 67.165 ;
        RECT 232.600 67.135 251.270 67.145 ;
        RECT 262.330 67.135 298.895 67.155 ;
        RECT 232.600 66.845 298.895 67.135 ;
        RECT 398.040 66.890 402.165 67.160 ;
        RECT 413.540 66.975 417.625 67.245 ;
        RECT 423.945 67.210 427.695 67.485 ;
        RECT 429.000 67.450 455.230 67.840 ;
        RECT 461.885 67.470 493.850 67.860 ;
        RECT 506.660 67.230 509.790 67.505 ;
        RECT 510.535 67.470 510.915 74.630 ;
        RECT 557.600 74.565 583.035 75.465 ;
        RECT 592.905 74.665 721.570 75.545 ;
        RECT 592.905 74.645 665.295 74.665 ;
        RECT 511.775 72.170 518.515 72.470 ;
        RECT 560.085 72.385 561.285 72.765 ;
        RECT 563.040 72.170 565.315 72.680 ;
        RECT 567.940 72.170 570.240 72.680 ;
        RECT 572.535 72.170 574.815 72.680 ;
        RECT 579.610 72.485 580.845 72.865 ;
        RECT 512.365 70.375 515.820 70.815 ;
        RECT 516.110 70.175 516.490 70.555 ;
        RECT 518.825 70.215 519.205 70.595 ;
        RECT 523.010 70.165 523.390 70.545 ;
        RECT 513.435 69.750 515.175 70.040 ;
        RECT 517.225 69.700 518.425 69.990 ;
        RECT 519.935 69.670 522.560 70.080 ;
        RECT 524.145 69.765 524.525 70.145 ;
        RECT 560.085 70.085 563.345 70.465 ;
        RECT 564.085 70.085 567.345 70.465 ;
        RECT 573.585 70.085 576.845 70.465 ;
        RECT 577.585 70.085 580.845 70.465 ;
        RECT 511.180 68.990 527.100 69.290 ;
        RECT 511.715 68.245 528.660 68.545 ;
        RECT 560.750 68.170 587.045 68.510 ;
        RECT 522.120 67.230 529.820 67.505 ;
        RECT 593.275 67.485 593.655 74.645 ;
        RECT 595.105 70.430 598.480 70.830 ;
        RECT 598.850 70.190 599.230 70.570 ;
        RECT 601.565 70.230 601.945 70.610 ;
        RECT 605.750 70.180 606.130 70.560 ;
        RECT 596.175 69.765 597.915 70.055 ;
        RECT 599.965 69.715 601.165 70.005 ;
        RECT 602.675 69.685 605.285 70.110 ;
        RECT 606.885 69.780 607.265 70.160 ;
        RECT 594.420 69.005 607.985 69.320 ;
        RECT 594.415 68.260 607.975 68.560 ;
        RECT 594.435 67.545 601.160 67.845 ;
        RECT 604.860 67.245 607.965 67.520 ;
        RECT 608.735 67.485 609.115 74.645 ;
        RECT 662.200 73.660 690.975 73.680 ;
        RECT 625.375 73.395 690.975 73.660 ;
        RECT 625.375 73.375 662.925 73.395 ;
        RECT 692.645 73.375 699.350 73.675 ;
        RECT 626.885 72.465 628.340 72.845 ;
        RECT 629.080 72.465 630.280 72.845 ;
        RECT 632.035 72.250 634.310 72.760 ;
        RECT 636.935 72.250 639.235 72.760 ;
        RECT 641.530 72.250 643.810 72.760 ;
        RECT 648.605 72.565 649.840 72.945 ;
        RECT 650.580 72.565 651.860 72.945 ;
        RECT 665.505 72.485 666.960 72.865 ;
        RECT 670.655 72.270 672.930 72.780 ;
        RECT 675.555 72.270 677.855 72.780 ;
        RECT 680.150 72.270 682.430 72.780 ;
        RECT 689.200 72.585 690.480 72.965 ;
        RECT 650.020 72.210 650.400 72.245 ;
        RECT 688.640 72.230 689.020 72.265 ;
        RECT 628.520 72.105 628.900 72.145 ;
        RECT 628.450 71.800 631.285 72.105 ;
        RECT 647.265 71.900 650.400 72.210 ;
        RECT 667.140 72.125 667.520 72.165 ;
        RECT 650.020 71.865 650.400 71.900 ;
        RECT 667.070 71.820 669.905 72.125 ;
        RECT 685.885 71.920 689.020 72.230 ;
        RECT 688.640 71.885 689.020 71.920 ;
        RECT 628.520 71.765 628.900 71.800 ;
        RECT 667.140 71.785 667.520 71.820 ;
        RECT 610.565 70.390 613.970 70.830 ;
        RECT 614.310 70.190 614.690 70.570 ;
        RECT 617.025 70.230 617.405 70.610 ;
        RECT 621.210 70.180 621.590 70.560 ;
        RECT 627.045 70.165 628.340 70.545 ;
        RECT 629.080 70.165 632.340 70.545 ;
        RECT 633.080 70.165 636.340 70.545 ;
        RECT 637.080 70.165 638.265 70.545 ;
        RECT 640.530 70.165 641.840 70.545 ;
        RECT 642.580 70.165 645.840 70.545 ;
        RECT 646.580 70.165 649.840 70.545 ;
        RECT 650.580 70.165 651.595 70.545 ;
        RECT 665.665 70.185 666.960 70.565 ;
        RECT 671.700 70.185 674.960 70.565 ;
        RECT 675.700 70.185 676.885 70.565 ;
        RECT 679.150 70.185 680.460 70.565 ;
        RECT 681.200 70.185 684.460 70.565 ;
        RECT 689.200 70.185 690.215 70.565 ;
        RECT 693.280 70.430 696.695 70.850 ;
        RECT 697.025 70.210 697.405 70.590 ;
        RECT 699.740 70.250 700.120 70.630 ;
        RECT 703.925 70.200 704.305 70.580 ;
        RECT 611.635 69.765 613.375 70.055 ;
        RECT 615.425 69.715 616.625 70.005 ;
        RECT 618.135 69.685 620.730 70.060 ;
        RECT 622.345 69.780 622.725 70.160 ;
        RECT 628.520 69.465 628.900 69.845 ;
        RECT 632.520 69.465 632.900 69.845 ;
        RECT 636.520 69.800 636.900 69.845 ;
        RECT 642.020 69.800 642.400 69.845 ;
        RECT 636.470 69.485 642.405 69.800 ;
        RECT 636.520 69.465 636.900 69.485 ;
        RECT 642.020 69.465 642.400 69.485 ;
        RECT 646.020 69.465 646.400 69.845 ;
        RECT 650.020 69.465 650.400 69.845 ;
        RECT 667.140 69.485 667.520 69.865 ;
        RECT 671.140 69.485 671.520 69.865 ;
        RECT 675.140 69.820 675.520 69.865 ;
        RECT 680.640 69.820 681.020 69.865 ;
        RECT 675.090 69.505 681.025 69.820 ;
        RECT 675.140 69.485 675.520 69.505 ;
        RECT 680.640 69.485 681.020 69.505 ;
        RECT 684.640 69.485 685.020 69.865 ;
        RECT 688.640 69.485 689.020 69.865 ;
        RECT 694.350 69.785 696.090 70.075 ;
        RECT 698.140 69.735 699.340 70.025 ;
        RECT 700.850 69.695 703.480 70.150 ;
        RECT 705.060 69.800 705.440 70.180 ;
        RECT 609.875 69.005 623.700 69.305 ;
        RECT 625.375 68.840 641.385 69.215 ;
        RECT 659.230 68.860 680.005 69.235 ;
        RECT 609.880 68.260 628.300 68.560 ;
        RECT 629.745 68.250 657.055 68.590 ;
        RECT 609.360 67.545 616.620 67.845 ;
        RECT 458.730 67.105 486.290 67.115 ;
        RECT 429.000 67.085 447.670 67.095 ;
        RECT 458.730 67.085 495.295 67.105 ;
        RECT 36.235 66.825 66.255 66.845 ;
        RECT 232.600 66.825 262.620 66.845 ;
        RECT 429.000 66.795 495.295 67.085 ;
        RECT 594.415 66.925 598.540 67.195 ;
        RECT 609.915 67.010 614.000 67.280 ;
        RECT 620.320 67.245 624.070 67.520 ;
        RECT 625.375 67.485 651.605 67.875 ;
        RECT 658.260 67.505 690.225 67.895 ;
        RECT 703.035 67.265 706.165 67.540 ;
        RECT 706.910 67.505 707.290 74.665 ;
        RECT 753.965 74.570 779.400 75.470 ;
        RECT 789.245 74.665 917.910 75.545 ;
        RECT 789.245 74.645 861.635 74.665 ;
        RECT 708.150 72.205 714.890 72.505 ;
        RECT 756.450 72.390 757.650 72.770 ;
        RECT 759.405 72.175 761.680 72.685 ;
        RECT 764.305 72.175 766.605 72.685 ;
        RECT 768.900 72.175 771.180 72.685 ;
        RECT 775.975 72.490 777.210 72.870 ;
        RECT 708.740 70.410 712.195 70.850 ;
        RECT 712.485 70.210 712.865 70.590 ;
        RECT 715.200 70.250 715.580 70.630 ;
        RECT 719.385 70.200 719.765 70.580 ;
        RECT 709.810 69.785 711.550 70.075 ;
        RECT 713.600 69.735 714.800 70.025 ;
        RECT 716.310 69.705 718.935 70.115 ;
        RECT 720.520 69.800 720.900 70.180 ;
        RECT 756.450 70.090 759.710 70.470 ;
        RECT 760.450 70.090 763.710 70.470 ;
        RECT 769.950 70.090 773.210 70.470 ;
        RECT 773.950 70.090 777.210 70.470 ;
        RECT 707.555 69.025 723.475 69.325 ;
        RECT 708.090 68.280 725.035 68.580 ;
        RECT 757.115 68.175 783.410 68.515 ;
        RECT 718.495 67.265 726.195 67.540 ;
        RECT 789.615 67.485 789.995 74.645 ;
        RECT 791.445 70.430 794.820 70.830 ;
        RECT 795.190 70.190 795.570 70.570 ;
        RECT 797.905 70.230 798.285 70.610 ;
        RECT 802.090 70.180 802.470 70.560 ;
        RECT 792.515 69.765 794.255 70.055 ;
        RECT 796.305 69.715 797.505 70.005 ;
        RECT 799.015 69.685 801.625 70.110 ;
        RECT 803.225 69.780 803.605 70.160 ;
        RECT 790.760 69.005 804.325 69.320 ;
        RECT 790.755 68.260 804.315 68.560 ;
        RECT 790.775 67.545 797.500 67.845 ;
        RECT 801.200 67.245 804.305 67.520 ;
        RECT 805.075 67.485 805.455 74.645 ;
        RECT 858.540 73.660 887.315 73.680 ;
        RECT 821.715 73.395 887.315 73.660 ;
        RECT 821.715 73.375 859.265 73.395 ;
        RECT 888.985 73.375 895.690 73.675 ;
        RECT 823.225 72.465 824.680 72.845 ;
        RECT 825.420 72.465 826.620 72.845 ;
        RECT 828.375 72.250 830.650 72.760 ;
        RECT 833.275 72.250 835.575 72.760 ;
        RECT 837.870 72.250 840.150 72.760 ;
        RECT 844.945 72.565 846.180 72.945 ;
        RECT 846.920 72.565 848.200 72.945 ;
        RECT 861.845 72.485 863.300 72.865 ;
        RECT 866.995 72.270 869.270 72.780 ;
        RECT 871.895 72.270 874.195 72.780 ;
        RECT 876.490 72.270 878.770 72.780 ;
        RECT 885.540 72.585 886.820 72.965 ;
        RECT 846.360 72.210 846.740 72.245 ;
        RECT 884.980 72.230 885.360 72.265 ;
        RECT 824.860 72.105 825.240 72.145 ;
        RECT 824.790 71.800 827.625 72.105 ;
        RECT 843.605 71.900 846.740 72.210 ;
        RECT 863.480 72.125 863.860 72.165 ;
        RECT 846.360 71.865 846.740 71.900 ;
        RECT 863.410 71.820 866.245 72.125 ;
        RECT 882.225 71.920 885.360 72.230 ;
        RECT 884.980 71.885 885.360 71.920 ;
        RECT 824.860 71.765 825.240 71.800 ;
        RECT 863.480 71.785 863.860 71.820 ;
        RECT 806.905 70.390 810.310 70.830 ;
        RECT 810.650 70.190 811.030 70.570 ;
        RECT 813.365 70.230 813.745 70.610 ;
        RECT 817.550 70.180 817.930 70.560 ;
        RECT 823.385 70.165 824.680 70.545 ;
        RECT 825.420 70.165 828.680 70.545 ;
        RECT 829.420 70.165 832.680 70.545 ;
        RECT 833.420 70.165 834.605 70.545 ;
        RECT 836.870 70.165 838.180 70.545 ;
        RECT 838.920 70.165 842.180 70.545 ;
        RECT 842.920 70.165 846.180 70.545 ;
        RECT 846.920 70.165 847.935 70.545 ;
        RECT 862.005 70.185 863.300 70.565 ;
        RECT 868.040 70.185 871.300 70.565 ;
        RECT 872.040 70.185 873.225 70.565 ;
        RECT 875.490 70.185 876.800 70.565 ;
        RECT 877.540 70.185 880.800 70.565 ;
        RECT 885.540 70.185 886.555 70.565 ;
        RECT 889.620 70.430 893.035 70.850 ;
        RECT 893.365 70.210 893.745 70.590 ;
        RECT 896.080 70.250 896.460 70.630 ;
        RECT 900.265 70.200 900.645 70.580 ;
        RECT 807.975 69.765 809.715 70.055 ;
        RECT 811.765 69.715 812.965 70.005 ;
        RECT 814.475 69.685 817.070 70.060 ;
        RECT 818.685 69.780 819.065 70.160 ;
        RECT 824.860 69.465 825.240 69.845 ;
        RECT 828.860 69.465 829.240 69.845 ;
        RECT 832.860 69.800 833.240 69.845 ;
        RECT 838.360 69.800 838.740 69.845 ;
        RECT 832.810 69.485 838.745 69.800 ;
        RECT 832.860 69.465 833.240 69.485 ;
        RECT 838.360 69.465 838.740 69.485 ;
        RECT 842.360 69.465 842.740 69.845 ;
        RECT 846.360 69.465 846.740 69.845 ;
        RECT 863.480 69.485 863.860 69.865 ;
        RECT 867.480 69.485 867.860 69.865 ;
        RECT 871.480 69.820 871.860 69.865 ;
        RECT 876.980 69.820 877.360 69.865 ;
        RECT 871.430 69.505 877.365 69.820 ;
        RECT 871.480 69.485 871.860 69.505 ;
        RECT 876.980 69.485 877.360 69.505 ;
        RECT 880.980 69.485 881.360 69.865 ;
        RECT 884.980 69.485 885.360 69.865 ;
        RECT 890.690 69.785 892.430 70.075 ;
        RECT 894.480 69.735 895.680 70.025 ;
        RECT 897.190 69.695 899.820 70.150 ;
        RECT 901.400 69.800 901.780 70.180 ;
        RECT 806.215 69.005 820.040 69.305 ;
        RECT 821.715 68.840 837.725 69.215 ;
        RECT 855.570 68.860 876.345 69.235 ;
        RECT 806.220 68.260 824.640 68.560 ;
        RECT 826.085 68.250 853.395 68.590 ;
        RECT 805.700 67.545 812.960 67.845 ;
        RECT 655.105 67.140 682.665 67.150 ;
        RECT 625.375 67.120 644.045 67.130 ;
        RECT 655.105 67.120 691.670 67.140 ;
        RECT 625.375 66.830 691.670 67.120 ;
        RECT 790.755 66.925 794.880 67.195 ;
        RECT 806.255 67.010 810.340 67.280 ;
        RECT 816.660 67.245 820.410 67.520 ;
        RECT 821.715 67.485 847.945 67.875 ;
        RECT 854.600 67.505 886.565 67.895 ;
        RECT 899.375 67.265 902.505 67.540 ;
        RECT 903.250 67.505 903.630 74.665 ;
        RECT 950.350 74.555 975.785 75.455 ;
        RECT 985.585 74.665 1114.250 75.545 ;
        RECT 985.585 74.645 1057.975 74.665 ;
        RECT 904.490 72.205 911.230 72.505 ;
        RECT 952.835 72.375 954.035 72.755 ;
        RECT 955.790 72.160 958.065 72.670 ;
        RECT 960.690 72.160 962.990 72.670 ;
        RECT 965.285 72.160 967.565 72.670 ;
        RECT 972.360 72.475 973.595 72.855 ;
        RECT 905.080 70.410 908.535 70.850 ;
        RECT 908.825 70.210 909.205 70.590 ;
        RECT 911.540 70.250 911.920 70.630 ;
        RECT 915.725 70.200 916.105 70.580 ;
        RECT 906.150 69.785 907.890 70.075 ;
        RECT 909.940 69.735 911.140 70.025 ;
        RECT 912.650 69.705 915.275 70.115 ;
        RECT 916.860 69.800 917.240 70.180 ;
        RECT 952.835 70.075 956.095 70.455 ;
        RECT 956.835 70.075 960.095 70.455 ;
        RECT 966.335 70.075 969.595 70.455 ;
        RECT 970.335 70.075 973.595 70.455 ;
        RECT 903.895 69.025 919.815 69.325 ;
        RECT 904.430 68.280 921.375 68.580 ;
        RECT 953.500 68.160 979.795 68.500 ;
        RECT 914.835 67.265 922.535 67.540 ;
        RECT 985.955 67.485 986.335 74.645 ;
        RECT 987.785 70.430 991.160 70.830 ;
        RECT 991.530 70.190 991.910 70.570 ;
        RECT 994.245 70.230 994.625 70.610 ;
        RECT 998.430 70.180 998.810 70.560 ;
        RECT 988.855 69.765 990.595 70.055 ;
        RECT 992.645 69.715 993.845 70.005 ;
        RECT 995.355 69.685 997.965 70.110 ;
        RECT 999.565 69.780 999.945 70.160 ;
        RECT 987.100 69.005 1000.665 69.320 ;
        RECT 987.095 68.260 1000.655 68.560 ;
        RECT 987.115 67.545 993.840 67.845 ;
        RECT 997.540 67.245 1000.645 67.520 ;
        RECT 1001.415 67.485 1001.795 74.645 ;
        RECT 1054.880 73.660 1083.655 73.680 ;
        RECT 1018.055 73.395 1083.655 73.660 ;
        RECT 1018.055 73.375 1055.605 73.395 ;
        RECT 1085.325 73.375 1092.030 73.675 ;
        RECT 1019.565 72.465 1021.020 72.845 ;
        RECT 1021.760 72.465 1022.960 72.845 ;
        RECT 1024.715 72.250 1026.990 72.760 ;
        RECT 1029.615 72.250 1031.915 72.760 ;
        RECT 1034.210 72.250 1036.490 72.760 ;
        RECT 1041.285 72.565 1042.520 72.945 ;
        RECT 1043.260 72.565 1044.540 72.945 ;
        RECT 1058.185 72.485 1059.640 72.865 ;
        RECT 1063.335 72.270 1065.610 72.780 ;
        RECT 1068.235 72.270 1070.535 72.780 ;
        RECT 1072.830 72.270 1075.110 72.780 ;
        RECT 1081.880 72.585 1083.160 72.965 ;
        RECT 1042.700 72.210 1043.080 72.245 ;
        RECT 1081.320 72.230 1081.700 72.265 ;
        RECT 1021.200 72.105 1021.580 72.145 ;
        RECT 1021.130 71.800 1023.965 72.105 ;
        RECT 1039.945 71.900 1043.080 72.210 ;
        RECT 1059.820 72.125 1060.200 72.165 ;
        RECT 1042.700 71.865 1043.080 71.900 ;
        RECT 1059.750 71.820 1062.585 72.125 ;
        RECT 1078.565 71.920 1081.700 72.230 ;
        RECT 1081.320 71.885 1081.700 71.920 ;
        RECT 1021.200 71.765 1021.580 71.800 ;
        RECT 1059.820 71.785 1060.200 71.820 ;
        RECT 1003.245 70.390 1006.650 70.830 ;
        RECT 1006.990 70.190 1007.370 70.570 ;
        RECT 1009.705 70.230 1010.085 70.610 ;
        RECT 1013.890 70.180 1014.270 70.560 ;
        RECT 1019.725 70.165 1021.020 70.545 ;
        RECT 1021.760 70.165 1025.020 70.545 ;
        RECT 1025.760 70.165 1029.020 70.545 ;
        RECT 1029.760 70.165 1030.945 70.545 ;
        RECT 1033.210 70.165 1034.520 70.545 ;
        RECT 1035.260 70.165 1038.520 70.545 ;
        RECT 1039.260 70.165 1042.520 70.545 ;
        RECT 1043.260 70.165 1044.275 70.545 ;
        RECT 1058.345 70.185 1059.640 70.565 ;
        RECT 1064.380 70.185 1067.640 70.565 ;
        RECT 1068.380 70.185 1069.565 70.565 ;
        RECT 1071.830 70.185 1073.140 70.565 ;
        RECT 1073.880 70.185 1077.140 70.565 ;
        RECT 1081.880 70.185 1082.895 70.565 ;
        RECT 1085.960 70.430 1089.375 70.850 ;
        RECT 1089.705 70.210 1090.085 70.590 ;
        RECT 1092.420 70.250 1092.800 70.630 ;
        RECT 1096.605 70.200 1096.985 70.580 ;
        RECT 1004.315 69.765 1006.055 70.055 ;
        RECT 1008.105 69.715 1009.305 70.005 ;
        RECT 1010.815 69.685 1013.410 70.060 ;
        RECT 1015.025 69.780 1015.405 70.160 ;
        RECT 1021.200 69.465 1021.580 69.845 ;
        RECT 1025.200 69.465 1025.580 69.845 ;
        RECT 1029.200 69.800 1029.580 69.845 ;
        RECT 1034.700 69.800 1035.080 69.845 ;
        RECT 1029.150 69.485 1035.085 69.800 ;
        RECT 1029.200 69.465 1029.580 69.485 ;
        RECT 1034.700 69.465 1035.080 69.485 ;
        RECT 1038.700 69.465 1039.080 69.845 ;
        RECT 1042.700 69.465 1043.080 69.845 ;
        RECT 1059.820 69.485 1060.200 69.865 ;
        RECT 1063.820 69.485 1064.200 69.865 ;
        RECT 1067.820 69.820 1068.200 69.865 ;
        RECT 1073.320 69.820 1073.700 69.865 ;
        RECT 1067.770 69.505 1073.705 69.820 ;
        RECT 1067.820 69.485 1068.200 69.505 ;
        RECT 1073.320 69.485 1073.700 69.505 ;
        RECT 1077.320 69.485 1077.700 69.865 ;
        RECT 1081.320 69.485 1081.700 69.865 ;
        RECT 1087.030 69.785 1088.770 70.075 ;
        RECT 1090.820 69.735 1092.020 70.025 ;
        RECT 1093.530 69.695 1096.160 70.150 ;
        RECT 1097.740 69.800 1098.120 70.180 ;
        RECT 1002.555 69.005 1016.380 69.305 ;
        RECT 1018.055 68.840 1034.065 69.215 ;
        RECT 1051.910 68.860 1072.685 69.235 ;
        RECT 1002.560 68.260 1020.980 68.560 ;
        RECT 1022.425 68.250 1049.735 68.590 ;
        RECT 1002.040 67.545 1009.300 67.845 ;
        RECT 851.445 67.140 879.005 67.150 ;
        RECT 821.715 67.120 840.385 67.130 ;
        RECT 851.445 67.120 888.010 67.140 ;
        RECT 821.715 66.830 888.010 67.120 ;
        RECT 987.095 66.925 991.220 67.195 ;
        RECT 1002.595 67.010 1006.680 67.280 ;
        RECT 1013.000 67.245 1016.750 67.520 ;
        RECT 1018.055 67.485 1044.285 67.875 ;
        RECT 1050.940 67.505 1082.905 67.895 ;
        RECT 1095.715 67.265 1098.845 67.540 ;
        RECT 1099.590 67.505 1099.970 74.665 ;
        RECT 1146.675 74.560 1172.110 75.460 ;
        RECT 1181.925 74.665 1310.590 75.545 ;
        RECT 1181.925 74.645 1254.315 74.665 ;
        RECT 1100.830 72.205 1107.570 72.505 ;
        RECT 1149.160 72.380 1150.360 72.760 ;
        RECT 1152.115 72.165 1154.390 72.675 ;
        RECT 1157.015 72.165 1159.315 72.675 ;
        RECT 1161.610 72.165 1163.890 72.675 ;
        RECT 1168.685 72.480 1169.920 72.860 ;
        RECT 1101.420 70.410 1104.875 70.850 ;
        RECT 1105.165 70.210 1105.545 70.590 ;
        RECT 1107.880 70.250 1108.260 70.630 ;
        RECT 1112.065 70.200 1112.445 70.580 ;
        RECT 1102.490 69.785 1104.230 70.075 ;
        RECT 1106.280 69.735 1107.480 70.025 ;
        RECT 1108.990 69.705 1111.615 70.115 ;
        RECT 1113.200 69.800 1113.580 70.180 ;
        RECT 1149.160 70.080 1152.420 70.460 ;
        RECT 1153.160 70.080 1156.420 70.460 ;
        RECT 1162.660 70.080 1165.920 70.460 ;
        RECT 1166.660 70.080 1169.920 70.460 ;
        RECT 1100.235 69.025 1116.155 69.325 ;
        RECT 1100.770 68.280 1117.715 68.580 ;
        RECT 1149.825 68.165 1176.120 68.505 ;
        RECT 1111.175 67.265 1118.875 67.540 ;
        RECT 1182.295 67.485 1182.675 74.645 ;
        RECT 1184.125 70.430 1187.500 70.830 ;
        RECT 1187.870 70.190 1188.250 70.570 ;
        RECT 1190.585 70.230 1190.965 70.610 ;
        RECT 1194.770 70.180 1195.150 70.560 ;
        RECT 1185.195 69.765 1186.935 70.055 ;
        RECT 1188.985 69.715 1190.185 70.005 ;
        RECT 1191.695 69.685 1194.305 70.110 ;
        RECT 1195.905 69.780 1196.285 70.160 ;
        RECT 1183.440 69.005 1197.005 69.320 ;
        RECT 1183.435 68.260 1196.995 68.560 ;
        RECT 1183.455 67.545 1190.180 67.845 ;
        RECT 1193.880 67.245 1196.985 67.520 ;
        RECT 1197.755 67.485 1198.135 74.645 ;
        RECT 1251.220 73.660 1279.995 73.680 ;
        RECT 1214.395 73.395 1279.995 73.660 ;
        RECT 1214.395 73.375 1251.945 73.395 ;
        RECT 1281.665 73.375 1288.370 73.675 ;
        RECT 1215.905 72.465 1217.360 72.845 ;
        RECT 1218.100 72.465 1219.300 72.845 ;
        RECT 1221.055 72.250 1223.330 72.760 ;
        RECT 1225.955 72.250 1228.255 72.760 ;
        RECT 1230.550 72.250 1232.830 72.760 ;
        RECT 1237.625 72.565 1238.860 72.945 ;
        RECT 1239.600 72.565 1240.880 72.945 ;
        RECT 1254.525 72.485 1255.980 72.865 ;
        RECT 1256.720 72.485 1257.920 72.865 ;
        RECT 1259.675 72.270 1261.950 72.780 ;
        RECT 1264.575 72.270 1266.875 72.780 ;
        RECT 1269.170 72.270 1271.450 72.780 ;
        RECT 1276.245 72.585 1277.480 72.965 ;
        RECT 1278.220 72.585 1279.500 72.965 ;
        RECT 1239.040 72.210 1239.420 72.245 ;
        RECT 1277.660 72.230 1278.040 72.265 ;
        RECT 1217.540 72.105 1217.920 72.145 ;
        RECT 1217.470 71.800 1220.305 72.105 ;
        RECT 1236.285 71.900 1239.420 72.210 ;
        RECT 1256.160 72.125 1256.540 72.165 ;
        RECT 1239.040 71.865 1239.420 71.900 ;
        RECT 1256.090 71.820 1258.925 72.125 ;
        RECT 1274.905 71.920 1278.040 72.230 ;
        RECT 1277.660 71.885 1278.040 71.920 ;
        RECT 1217.540 71.765 1217.920 71.800 ;
        RECT 1256.160 71.785 1256.540 71.820 ;
        RECT 1199.585 70.390 1202.990 70.830 ;
        RECT 1203.330 70.190 1203.710 70.570 ;
        RECT 1206.045 70.230 1206.425 70.610 ;
        RECT 1210.230 70.180 1210.610 70.560 ;
        RECT 1216.065 70.165 1217.360 70.545 ;
        RECT 1218.100 70.165 1221.360 70.545 ;
        RECT 1222.100 70.165 1225.360 70.545 ;
        RECT 1226.100 70.165 1227.285 70.545 ;
        RECT 1229.550 70.165 1230.860 70.545 ;
        RECT 1231.600 70.165 1234.860 70.545 ;
        RECT 1235.600 70.165 1238.860 70.545 ;
        RECT 1239.600 70.165 1240.615 70.545 ;
        RECT 1254.685 70.185 1255.980 70.565 ;
        RECT 1256.720 70.185 1259.980 70.565 ;
        RECT 1260.720 70.185 1263.980 70.565 ;
        RECT 1264.720 70.185 1265.905 70.565 ;
        RECT 1268.170 70.185 1269.480 70.565 ;
        RECT 1270.220 70.185 1273.480 70.565 ;
        RECT 1274.220 70.185 1277.480 70.565 ;
        RECT 1278.220 70.185 1279.235 70.565 ;
        RECT 1282.300 70.430 1285.715 70.850 ;
        RECT 1286.045 70.210 1286.425 70.590 ;
        RECT 1288.760 70.250 1289.140 70.630 ;
        RECT 1292.945 70.200 1293.325 70.580 ;
        RECT 1200.655 69.765 1202.395 70.055 ;
        RECT 1204.445 69.715 1205.645 70.005 ;
        RECT 1207.155 69.685 1209.750 70.060 ;
        RECT 1211.365 69.780 1211.745 70.160 ;
        RECT 1217.540 69.465 1217.920 69.845 ;
        RECT 1221.540 69.465 1221.920 69.845 ;
        RECT 1225.540 69.800 1225.920 69.845 ;
        RECT 1231.040 69.800 1231.420 69.845 ;
        RECT 1225.490 69.485 1231.425 69.800 ;
        RECT 1225.540 69.465 1225.920 69.485 ;
        RECT 1231.040 69.465 1231.420 69.485 ;
        RECT 1235.040 69.465 1235.420 69.845 ;
        RECT 1239.040 69.465 1239.420 69.845 ;
        RECT 1256.160 69.485 1256.540 69.865 ;
        RECT 1260.160 69.485 1260.540 69.865 ;
        RECT 1264.160 69.820 1264.540 69.865 ;
        RECT 1269.660 69.820 1270.040 69.865 ;
        RECT 1264.110 69.505 1270.045 69.820 ;
        RECT 1264.160 69.485 1264.540 69.505 ;
        RECT 1269.660 69.485 1270.040 69.505 ;
        RECT 1273.660 69.485 1274.040 69.865 ;
        RECT 1277.660 69.485 1278.040 69.865 ;
        RECT 1283.370 69.785 1285.110 70.075 ;
        RECT 1287.160 69.735 1288.360 70.025 ;
        RECT 1289.870 69.695 1292.500 70.150 ;
        RECT 1294.080 69.800 1294.460 70.180 ;
        RECT 1198.895 69.005 1212.720 69.305 ;
        RECT 1214.395 68.840 1230.405 69.215 ;
        RECT 1248.250 68.860 1269.025 69.235 ;
        RECT 1281.650 69.025 1295.265 69.325 ;
        RECT 1198.900 68.260 1217.320 68.560 ;
        RECT 1218.765 68.250 1246.075 68.590 ;
        RECT 1257.385 68.270 1279.940 68.610 ;
        RECT 1281.050 68.280 1295.695 68.580 ;
        RECT 1198.380 67.545 1205.640 67.845 ;
        RECT 1047.785 67.140 1075.345 67.150 ;
        RECT 1018.055 67.120 1036.725 67.130 ;
        RECT 1047.785 67.120 1084.350 67.140 ;
        RECT 1018.055 66.830 1084.350 67.120 ;
        RECT 1183.435 66.925 1187.560 67.195 ;
        RECT 1198.935 67.010 1203.020 67.280 ;
        RECT 1209.340 67.245 1213.090 67.520 ;
        RECT 1214.395 67.485 1240.625 67.875 ;
        RECT 1247.280 67.505 1279.245 67.895 ;
        RECT 1292.055 67.265 1295.185 67.540 ;
        RECT 1295.930 67.505 1296.310 74.665 ;
        RECT 1297.170 72.205 1303.910 72.505 ;
        RECT 1297.760 70.410 1301.215 70.850 ;
        RECT 1304.220 70.250 1304.600 70.630 ;
        RECT 1302.620 69.735 1303.820 70.025 ;
        RECT 1309.540 69.800 1309.920 70.180 ;
        RECT 1296.575 69.025 1312.495 69.325 ;
        RECT 1297.110 68.280 1314.055 68.580 ;
        RECT 1244.125 67.140 1271.685 67.150 ;
        RECT 1214.395 67.120 1233.065 67.130 ;
        RECT 1244.125 67.120 1280.690 67.140 ;
        RECT 1214.395 66.830 1280.690 67.120 ;
        RECT 625.375 66.810 655.395 66.830 ;
        RECT 821.715 66.810 851.735 66.830 ;
        RECT 1018.055 66.810 1048.075 66.830 ;
        RECT 1214.395 66.810 1244.415 66.830 ;
        RECT 429.000 66.775 459.020 66.795 ;
        RECT 6.510 66.365 10.640 66.665 ;
        RECT -59.735 65.455 -56.170 65.465 ;
        RECT -59.735 65.130 -55.375 65.455 ;
        RECT -9.410 65.210 -3.495 65.545 ;
        RECT -6.140 65.190 -3.495 65.210 ;
        RECT -56.330 65.120 -55.375 65.130 ;
        RECT -79.140 64.490 -75.840 64.870 ;
        RECT -75.140 64.490 -71.840 64.870 ;
        RECT -65.640 64.490 -62.340 64.870 ;
        RECT -61.640 64.490 -58.340 64.870 ;
        RECT -28.815 64.570 -25.515 64.950 ;
        RECT -24.815 64.570 -21.515 64.950 ;
        RECT -15.315 64.570 -12.015 64.950 ;
        RECT -11.315 64.570 -8.015 64.950 ;
        RECT -79.140 62.490 -77.855 62.870 ;
        RECT -59.825 62.490 -58.340 62.870 ;
        RECT -28.815 62.570 -27.530 62.950 ;
        RECT -9.500 62.570 -8.015 62.950 ;
        RECT -77.635 61.810 -76.115 62.170 ;
        RECT -27.310 61.890 -25.790 62.250 ;
        RECT 4.135 60.535 4.515 66.365 ;
        RECT 13.015 66.315 17.515 66.625 ;
        RECT 21.970 66.365 26.100 66.665 ;
        RECT 8.975 65.765 15.365 66.055 ;
        RECT 8.390 65.185 19.045 65.520 ;
        RECT 7.740 64.600 10.660 64.900 ;
        RECT 14.205 64.585 17.575 64.885 ;
        RECT 5.955 63.850 6.335 64.230 ;
        RECT 8.360 63.865 10.140 64.155 ;
        RECT 11.615 63.955 12.805 64.240 ;
        RECT 15.735 63.835 17.045 64.155 ;
        RECT 7.090 63.250 7.470 63.630 ;
        RECT 10.835 63.290 11.215 63.670 ;
        RECT 13.545 63.280 13.925 63.660 ;
        RECT 14.955 63.125 18.135 63.445 ;
        RECT 4.885 60.535 8.980 60.540 ;
        RECT 19.595 60.535 19.975 66.365 ;
        RECT 28.475 66.315 32.975 66.625 ;
        RECT 120.145 66.385 124.275 66.685 ;
        RECT 71.185 66.155 102.930 66.175 ;
        RECT 24.435 65.765 30.825 66.055 ;
        RECT 35.705 65.905 102.930 66.155 ;
        RECT 35.705 65.885 71.615 65.905 ;
        RECT 107.150 65.785 113.540 66.075 ;
        RECT 23.850 65.185 34.355 65.520 ;
        RECT 59.325 65.320 69.875 65.655 ;
        RECT 106.565 65.205 117.045 65.540 ;
        RECT 23.200 64.600 26.120 64.900 ;
        RECT 29.665 64.585 33.035 64.885 ;
        RECT 37.915 64.680 39.220 65.060 ;
        RECT 39.920 64.680 43.220 65.060 ;
        RECT 43.920 64.680 47.220 65.060 ;
        RECT 47.920 64.680 49.280 65.060 ;
        RECT 51.255 64.680 52.720 65.060 ;
        RECT 53.420 64.680 56.720 65.060 ;
        RECT 57.420 64.680 60.720 65.060 ;
        RECT 61.420 64.680 62.600 65.060 ;
        RECT 76.535 64.700 77.840 65.080 ;
        RECT 82.540 64.700 85.840 65.080 ;
        RECT 86.540 64.700 87.900 65.080 ;
        RECT 89.875 64.700 91.340 65.080 ;
        RECT 92.040 64.700 95.340 65.080 ;
        RECT 100.040 64.700 101.220 65.080 ;
        RECT 39.380 64.335 39.760 64.370 ;
        RECT 21.415 63.850 21.795 64.230 ;
        RECT 23.820 63.865 25.600 64.155 ;
        RECT 27.075 63.955 28.265 64.240 ;
        RECT 31.195 63.835 32.505 64.155 ;
        RECT 39.115 64.025 42.125 64.335 ;
        RECT 39.380 63.990 39.760 64.025 ;
        RECT 43.380 63.990 44.470 64.370 ;
        RECT 47.380 64.365 47.760 64.370 ;
        RECT 44.900 64.000 47.765 64.365 ;
        RECT 52.880 64.345 53.260 64.370 ;
        RECT 52.865 64.025 55.010 64.345 ;
        RECT 47.380 63.990 47.760 64.000 ;
        RECT 52.880 63.990 53.260 64.025 ;
        RECT 55.925 63.990 57.260 64.370 ;
        RECT 60.880 64.350 61.260 64.370 ;
        RECT 78.000 64.355 78.380 64.390 ;
        RECT 58.415 64.030 61.325 64.350 ;
        RECT 77.735 64.045 80.745 64.355 ;
        RECT 60.880 63.990 61.260 64.030 ;
        RECT 78.000 64.010 78.380 64.045 ;
        RECT 82.000 64.010 83.090 64.390 ;
        RECT 86.000 64.385 86.380 64.390 ;
        RECT 83.520 64.020 86.385 64.385 ;
        RECT 91.500 64.365 91.880 64.390 ;
        RECT 91.485 64.045 93.630 64.365 ;
        RECT 86.000 64.010 86.380 64.020 ;
        RECT 91.500 64.010 91.880 64.045 ;
        RECT 94.545 64.010 95.880 64.390 ;
        RECT 99.500 64.370 99.880 64.390 ;
        RECT 97.035 64.050 99.945 64.370 ;
        RECT 99.500 64.010 99.880 64.050 ;
        RECT 104.130 63.870 104.510 64.250 ;
        RECT 106.535 63.885 108.315 64.175 ;
        RECT 109.790 63.975 110.980 64.260 ;
        RECT 113.910 63.855 115.220 64.175 ;
        RECT 22.550 63.250 22.930 63.630 ;
        RECT 26.295 63.290 26.675 63.670 ;
        RECT 29.005 63.280 29.385 63.660 ;
        RECT 30.415 63.125 33.595 63.445 ;
        RECT 105.265 63.270 105.645 63.650 ;
        RECT 109.010 63.310 109.390 63.690 ;
        RECT 111.720 63.300 112.100 63.680 ;
        RECT 113.130 63.145 116.310 63.465 ;
        RECT 37.730 62.680 39.220 63.060 ;
        RECT 39.920 62.680 41.205 63.060 ;
        RECT 59.235 62.680 60.720 63.060 ;
        RECT 61.420 62.680 62.495 63.060 ;
        RECT 76.350 62.700 77.840 63.080 ;
        RECT 100.040 62.700 101.115 63.080 ;
        RECT 39.380 61.990 40.470 62.370 ;
        RECT 41.425 62.000 42.945 62.360 ;
        RECT 43.865 61.995 56.715 62.330 ;
        RECT 60.880 62.325 61.260 62.370 ;
        RECT 60.145 62.025 61.455 62.325 ;
        RECT 60.880 61.990 61.260 62.025 ;
        RECT 78.000 62.010 79.090 62.390 ;
        RECT 80.045 62.020 81.565 62.380 ;
        RECT 82.485 62.015 95.335 62.350 ;
        RECT 99.500 62.345 99.880 62.390 ;
        RECT 98.765 62.045 100.075 62.345 ;
        RECT 99.500 62.010 99.880 62.045 ;
        RECT 68.560 61.480 101.510 61.515 ;
        RECT 36.235 61.150 101.510 61.480 ;
        RECT 36.235 61.130 69.315 61.150 ;
        RECT 103.305 61.140 107.565 61.495 ;
        RECT 101.510 60.555 107.155 60.560 ;
        RECT 117.770 60.555 118.150 66.385 ;
        RECT 126.650 66.335 131.150 66.645 ;
        RECT 202.875 66.365 207.005 66.665 ;
        RECT 122.610 65.785 129.000 66.075 ;
        RECT 122.025 65.205 138.045 65.540 ;
        RECT 186.760 65.220 192.675 65.555 ;
        RECT 190.030 65.200 192.675 65.220 ;
        RECT 121.375 64.620 124.295 64.920 ;
        RECT 127.840 64.605 131.210 64.905 ;
        RECT 167.355 64.580 170.655 64.960 ;
        RECT 171.355 64.580 174.655 64.960 ;
        RECT 180.855 64.580 184.155 64.960 ;
        RECT 184.855 64.580 188.155 64.960 ;
        RECT 119.590 63.870 119.970 64.250 ;
        RECT 121.995 63.885 123.775 64.175 ;
        RECT 125.250 63.975 126.440 64.260 ;
        RECT 129.370 63.855 130.680 64.175 ;
        RECT 120.725 63.270 121.105 63.650 ;
        RECT 124.470 63.310 124.850 63.690 ;
        RECT 127.180 63.300 127.560 63.680 ;
        RECT 128.590 63.145 131.770 63.465 ;
        RECT 167.355 62.580 168.640 62.960 ;
        RECT 186.670 62.580 188.155 62.960 ;
        RECT 118.870 62.060 123.020 62.330 ;
        RECT 168.860 61.900 170.380 62.260 ;
        RECT 118.520 60.555 122.615 60.560 ;
        RECT 74.855 60.550 107.155 60.555 ;
        RECT 117.400 60.550 122.615 60.555 ;
        RECT 20.345 60.535 24.440 60.540 ;
        RECT 74.855 60.535 132.430 60.550 ;
        RECT 200.500 60.535 200.880 66.365 ;
        RECT 209.380 66.315 213.880 66.625 ;
        RECT 218.335 66.365 222.465 66.665 ;
        RECT 205.340 65.765 211.730 66.055 ;
        RECT 204.755 65.185 215.410 65.520 ;
        RECT 204.105 64.600 207.025 64.900 ;
        RECT 210.570 64.585 213.940 64.885 ;
        RECT 202.320 63.850 202.700 64.230 ;
        RECT 204.725 63.865 206.505 64.155 ;
        RECT 207.980 63.955 209.170 64.240 ;
        RECT 212.100 63.835 213.410 64.155 ;
        RECT 203.455 63.250 203.835 63.630 ;
        RECT 207.200 63.290 207.580 63.670 ;
        RECT 209.910 63.280 210.290 63.660 ;
        RECT 211.320 63.125 214.500 63.445 ;
        RECT 201.250 60.535 205.345 60.540 ;
        RECT 215.960 60.535 216.340 66.365 ;
        RECT 224.840 66.315 229.340 66.625 ;
        RECT 316.510 66.385 320.640 66.685 ;
        RECT 267.550 66.155 299.295 66.175 ;
        RECT 220.800 65.765 227.190 66.055 ;
        RECT 232.070 65.905 299.295 66.155 ;
        RECT 232.070 65.885 267.980 65.905 ;
        RECT 303.515 65.785 309.905 66.075 ;
        RECT 220.215 65.185 230.720 65.520 ;
        RECT 255.690 65.320 266.240 65.655 ;
        RECT 302.930 65.205 313.410 65.540 ;
        RECT 219.565 64.600 222.485 64.900 ;
        RECT 226.030 64.585 229.400 64.885 ;
        RECT 234.280 64.680 235.585 65.060 ;
        RECT 236.285 64.680 239.585 65.060 ;
        RECT 240.285 64.680 243.585 65.060 ;
        RECT 244.285 64.680 245.645 65.060 ;
        RECT 247.620 64.680 249.085 65.060 ;
        RECT 249.785 64.680 253.085 65.060 ;
        RECT 253.785 64.680 257.085 65.060 ;
        RECT 257.785 64.680 258.965 65.060 ;
        RECT 272.900 64.700 274.205 65.080 ;
        RECT 278.905 64.700 282.205 65.080 ;
        RECT 282.905 64.700 284.265 65.080 ;
        RECT 286.240 64.700 287.705 65.080 ;
        RECT 288.405 64.700 291.705 65.080 ;
        RECT 296.405 64.700 297.585 65.080 ;
        RECT 235.745 64.335 236.125 64.370 ;
        RECT 217.780 63.850 218.160 64.230 ;
        RECT 220.185 63.865 221.965 64.155 ;
        RECT 223.440 63.955 224.630 64.240 ;
        RECT 227.560 63.835 228.870 64.155 ;
        RECT 235.480 64.025 238.490 64.335 ;
        RECT 235.745 63.990 236.125 64.025 ;
        RECT 239.745 63.990 240.835 64.370 ;
        RECT 243.745 64.365 244.125 64.370 ;
        RECT 241.265 64.000 244.130 64.365 ;
        RECT 249.245 64.345 249.625 64.370 ;
        RECT 249.230 64.025 251.375 64.345 ;
        RECT 243.745 63.990 244.125 64.000 ;
        RECT 249.245 63.990 249.625 64.025 ;
        RECT 252.290 63.990 253.625 64.370 ;
        RECT 257.245 64.350 257.625 64.370 ;
        RECT 274.365 64.355 274.745 64.390 ;
        RECT 254.780 64.030 257.690 64.350 ;
        RECT 274.100 64.045 277.110 64.355 ;
        RECT 257.245 63.990 257.625 64.030 ;
        RECT 274.365 64.010 274.745 64.045 ;
        RECT 278.365 64.010 279.455 64.390 ;
        RECT 282.365 64.385 282.745 64.390 ;
        RECT 279.885 64.020 282.750 64.385 ;
        RECT 287.865 64.365 288.245 64.390 ;
        RECT 287.850 64.045 289.995 64.365 ;
        RECT 282.365 64.010 282.745 64.020 ;
        RECT 287.865 64.010 288.245 64.045 ;
        RECT 290.910 64.010 292.245 64.390 ;
        RECT 295.865 64.370 296.245 64.390 ;
        RECT 293.400 64.050 296.310 64.370 ;
        RECT 295.865 64.010 296.245 64.050 ;
        RECT 300.495 63.870 300.875 64.250 ;
        RECT 302.900 63.885 304.680 64.175 ;
        RECT 306.155 63.975 307.345 64.260 ;
        RECT 310.275 63.855 311.585 64.175 ;
        RECT 218.915 63.250 219.295 63.630 ;
        RECT 222.660 63.290 223.040 63.670 ;
        RECT 225.370 63.280 225.750 63.660 ;
        RECT 226.780 63.125 229.960 63.445 ;
        RECT 301.630 63.270 302.010 63.650 ;
        RECT 305.375 63.310 305.755 63.690 ;
        RECT 308.085 63.300 308.465 63.680 ;
        RECT 309.495 63.145 312.675 63.465 ;
        RECT 234.095 62.680 235.585 63.060 ;
        RECT 236.285 62.680 237.570 63.060 ;
        RECT 255.600 62.680 257.085 63.060 ;
        RECT 257.785 62.680 258.860 63.060 ;
        RECT 272.715 62.700 274.205 63.080 ;
        RECT 296.405 62.700 297.480 63.080 ;
        RECT 235.745 61.990 236.835 62.370 ;
        RECT 237.790 62.000 239.310 62.360 ;
        RECT 240.230 61.995 253.080 62.330 ;
        RECT 257.245 62.325 257.625 62.370 ;
        RECT 256.510 62.025 257.820 62.325 ;
        RECT 257.245 61.990 257.625 62.025 ;
        RECT 274.365 62.010 275.455 62.390 ;
        RECT 276.410 62.020 277.930 62.380 ;
        RECT 278.850 62.015 291.700 62.350 ;
        RECT 295.865 62.345 296.245 62.390 ;
        RECT 295.130 62.045 296.440 62.345 ;
        RECT 295.865 62.010 296.245 62.045 ;
        RECT 264.925 61.480 297.875 61.515 ;
        RECT 232.600 61.150 297.875 61.480 ;
        RECT 232.600 61.130 265.680 61.150 ;
        RECT 299.670 61.140 303.930 61.495 ;
        RECT 297.875 60.555 303.520 60.560 ;
        RECT 314.135 60.555 314.515 66.385 ;
        RECT 323.015 66.335 327.515 66.645 ;
        RECT 399.275 66.315 403.405 66.615 ;
        RECT 318.975 65.785 325.365 66.075 ;
        RECT 318.390 65.205 334.410 65.540 ;
        RECT 383.150 65.180 389.065 65.515 ;
        RECT 386.420 65.160 389.065 65.180 ;
        RECT 317.740 64.620 320.660 64.920 ;
        RECT 324.205 64.605 327.575 64.905 ;
        RECT 363.745 64.540 367.045 64.920 ;
        RECT 367.745 64.540 371.045 64.920 ;
        RECT 377.245 64.540 380.545 64.920 ;
        RECT 381.245 64.540 384.545 64.920 ;
        RECT 315.955 63.870 316.335 64.250 ;
        RECT 318.360 63.885 320.140 64.175 ;
        RECT 321.615 63.975 322.805 64.260 ;
        RECT 325.735 63.855 327.045 64.175 ;
        RECT 317.090 63.270 317.470 63.650 ;
        RECT 320.835 63.310 321.215 63.690 ;
        RECT 323.545 63.300 323.925 63.680 ;
        RECT 324.955 63.145 328.135 63.465 ;
        RECT 363.745 62.540 365.030 62.920 ;
        RECT 383.060 62.540 384.545 62.920 ;
        RECT 315.235 62.060 319.385 62.330 ;
        RECT 365.250 61.860 366.770 62.220 ;
        RECT 314.885 60.555 318.980 60.560 ;
        RECT 271.220 60.550 303.520 60.555 ;
        RECT 313.765 60.550 318.980 60.555 ;
        RECT 216.710 60.535 220.805 60.540 ;
        RECT 271.220 60.535 328.795 60.550 ;
        RECT 3.765 60.530 8.980 60.535 ;
        RECT 19.225 60.530 24.440 60.535 ;
        RECT 34.685 60.530 132.430 60.535 ;
        RECT -82.825 59.445 -56.170 60.345 ;
        RECT -32.500 59.525 -5.845 60.425 ;
        RECT 3.765 59.655 132.430 60.530 ;
        RECT 200.130 60.530 205.345 60.535 ;
        RECT 215.590 60.530 220.805 60.535 ;
        RECT 231.050 60.530 328.795 60.535 ;
        RECT 3.765 59.635 74.935 59.655 ;
        RECT 163.670 59.535 190.325 60.435 ;
        RECT 200.130 59.655 328.795 60.530 ;
        RECT 396.900 60.485 397.280 66.315 ;
        RECT 405.780 66.265 410.280 66.575 ;
        RECT 414.735 66.315 418.865 66.615 ;
        RECT 401.740 65.715 408.130 66.005 ;
        RECT 401.155 65.135 411.810 65.470 ;
        RECT 400.505 64.550 403.425 64.850 ;
        RECT 406.970 64.535 410.340 64.835 ;
        RECT 398.720 63.800 399.100 64.180 ;
        RECT 401.125 63.815 402.905 64.105 ;
        RECT 404.380 63.905 405.570 64.190 ;
        RECT 408.500 63.785 409.810 64.105 ;
        RECT 399.855 63.200 400.235 63.580 ;
        RECT 403.600 63.240 403.980 63.620 ;
        RECT 406.310 63.230 406.690 63.610 ;
        RECT 407.720 63.075 410.900 63.395 ;
        RECT 397.650 60.485 401.745 60.490 ;
        RECT 412.360 60.485 412.740 66.315 ;
        RECT 421.240 66.265 425.740 66.575 ;
        RECT 512.910 66.335 517.040 66.635 ;
        RECT 463.950 66.105 495.695 66.125 ;
        RECT 417.200 65.715 423.590 66.005 ;
        RECT 428.470 65.855 495.695 66.105 ;
        RECT 428.470 65.835 464.380 65.855 ;
        RECT 499.915 65.735 506.305 66.025 ;
        RECT 416.615 65.135 427.120 65.470 ;
        RECT 452.090 65.270 462.640 65.605 ;
        RECT 499.330 65.155 509.810 65.490 ;
        RECT 415.965 64.550 418.885 64.850 ;
        RECT 422.430 64.535 425.800 64.835 ;
        RECT 430.680 64.630 431.985 65.010 ;
        RECT 432.685 64.630 435.985 65.010 ;
        RECT 436.685 64.630 439.985 65.010 ;
        RECT 440.685 64.630 442.045 65.010 ;
        RECT 444.020 64.630 445.485 65.010 ;
        RECT 446.185 64.630 449.485 65.010 ;
        RECT 450.185 64.630 453.485 65.010 ;
        RECT 454.185 64.630 455.365 65.010 ;
        RECT 469.300 64.650 470.605 65.030 ;
        RECT 475.305 64.650 478.605 65.030 ;
        RECT 479.305 64.650 480.665 65.030 ;
        RECT 482.640 64.650 484.105 65.030 ;
        RECT 484.805 64.650 488.105 65.030 ;
        RECT 492.805 64.650 493.985 65.030 ;
        RECT 432.145 64.285 432.525 64.320 ;
        RECT 414.180 63.800 414.560 64.180 ;
        RECT 416.585 63.815 418.365 64.105 ;
        RECT 419.840 63.905 421.030 64.190 ;
        RECT 423.960 63.785 425.270 64.105 ;
        RECT 431.880 63.975 434.890 64.285 ;
        RECT 432.145 63.940 432.525 63.975 ;
        RECT 436.145 63.940 437.235 64.320 ;
        RECT 440.145 64.315 440.525 64.320 ;
        RECT 437.665 63.950 440.530 64.315 ;
        RECT 445.645 64.295 446.025 64.320 ;
        RECT 445.630 63.975 447.775 64.295 ;
        RECT 440.145 63.940 440.525 63.950 ;
        RECT 445.645 63.940 446.025 63.975 ;
        RECT 448.690 63.940 450.025 64.320 ;
        RECT 453.645 64.300 454.025 64.320 ;
        RECT 470.765 64.305 471.145 64.340 ;
        RECT 451.180 63.980 454.090 64.300 ;
        RECT 470.500 63.995 473.510 64.305 ;
        RECT 453.645 63.940 454.025 63.980 ;
        RECT 470.765 63.960 471.145 63.995 ;
        RECT 474.765 63.960 475.855 64.340 ;
        RECT 478.765 64.335 479.145 64.340 ;
        RECT 476.285 63.970 479.150 64.335 ;
        RECT 484.265 64.315 484.645 64.340 ;
        RECT 484.250 63.995 486.395 64.315 ;
        RECT 478.765 63.960 479.145 63.970 ;
        RECT 484.265 63.960 484.645 63.995 ;
        RECT 487.310 63.960 488.645 64.340 ;
        RECT 492.265 64.320 492.645 64.340 ;
        RECT 489.800 64.000 492.710 64.320 ;
        RECT 492.265 63.960 492.645 64.000 ;
        RECT 496.895 63.820 497.275 64.200 ;
        RECT 499.300 63.835 501.080 64.125 ;
        RECT 502.555 63.925 503.745 64.210 ;
        RECT 506.675 63.805 507.985 64.125 ;
        RECT 415.315 63.200 415.695 63.580 ;
        RECT 419.060 63.240 419.440 63.620 ;
        RECT 421.770 63.230 422.150 63.610 ;
        RECT 423.180 63.075 426.360 63.395 ;
        RECT 498.030 63.220 498.410 63.600 ;
        RECT 501.775 63.260 502.155 63.640 ;
        RECT 504.485 63.250 504.865 63.630 ;
        RECT 505.895 63.095 509.075 63.415 ;
        RECT 430.495 62.630 431.985 63.010 ;
        RECT 432.685 62.630 433.970 63.010 ;
        RECT 452.000 62.630 453.485 63.010 ;
        RECT 454.185 62.630 455.260 63.010 ;
        RECT 469.115 62.650 470.605 63.030 ;
        RECT 492.805 62.650 493.880 63.030 ;
        RECT 432.145 61.940 433.235 62.320 ;
        RECT 434.190 61.950 435.710 62.310 ;
        RECT 436.630 61.945 449.480 62.280 ;
        RECT 453.645 62.275 454.025 62.320 ;
        RECT 452.910 61.975 454.220 62.275 ;
        RECT 453.645 61.940 454.025 61.975 ;
        RECT 470.765 61.960 471.855 62.340 ;
        RECT 472.810 61.970 474.330 62.330 ;
        RECT 475.250 61.965 488.100 62.300 ;
        RECT 492.265 62.295 492.645 62.340 ;
        RECT 491.530 61.995 492.840 62.295 ;
        RECT 492.265 61.960 492.645 61.995 ;
        RECT 461.325 61.430 494.275 61.465 ;
        RECT 429.000 61.100 494.275 61.430 ;
        RECT 429.000 61.080 462.080 61.100 ;
        RECT 496.070 61.090 500.330 61.445 ;
        RECT 494.275 60.505 499.920 60.510 ;
        RECT 510.535 60.505 510.915 66.335 ;
        RECT 519.415 66.285 523.915 66.595 ;
        RECT 595.650 66.350 599.780 66.650 ;
        RECT 515.375 65.735 521.765 66.025 ;
        RECT 514.790 65.155 530.810 65.490 ;
        RECT 579.470 65.225 585.385 65.560 ;
        RECT 582.740 65.205 585.385 65.225 ;
        RECT 514.140 64.570 517.060 64.870 ;
        RECT 520.605 64.555 523.975 64.855 ;
        RECT 560.065 64.585 563.365 64.965 ;
        RECT 564.065 64.585 567.365 64.965 ;
        RECT 573.565 64.585 576.865 64.965 ;
        RECT 577.565 64.585 580.865 64.965 ;
        RECT 512.355 63.820 512.735 64.200 ;
        RECT 514.760 63.835 516.540 64.125 ;
        RECT 518.015 63.925 519.205 64.210 ;
        RECT 522.135 63.805 523.445 64.125 ;
        RECT 513.490 63.220 513.870 63.600 ;
        RECT 517.235 63.260 517.615 63.640 ;
        RECT 519.945 63.250 520.325 63.630 ;
        RECT 521.355 63.095 524.535 63.415 ;
        RECT 560.065 62.585 561.350 62.965 ;
        RECT 579.380 62.585 580.865 62.965 ;
        RECT 511.635 62.010 515.785 62.280 ;
        RECT 561.570 61.905 563.090 62.265 ;
        RECT 593.275 60.520 593.655 66.350 ;
        RECT 602.155 66.300 606.655 66.610 ;
        RECT 611.110 66.350 615.240 66.650 ;
        RECT 598.115 65.750 604.505 66.040 ;
        RECT 597.530 65.170 608.185 65.505 ;
        RECT 596.880 64.585 599.800 64.885 ;
        RECT 603.345 64.570 606.715 64.870 ;
        RECT 595.095 63.835 595.475 64.215 ;
        RECT 597.500 63.850 599.280 64.140 ;
        RECT 600.755 63.940 601.945 64.225 ;
        RECT 604.875 63.820 606.185 64.140 ;
        RECT 596.230 63.235 596.610 63.615 ;
        RECT 599.975 63.275 600.355 63.655 ;
        RECT 602.685 63.265 603.065 63.645 ;
        RECT 604.095 63.110 607.275 63.430 ;
        RECT 594.025 60.520 598.120 60.525 ;
        RECT 608.735 60.520 609.115 66.350 ;
        RECT 617.615 66.300 622.115 66.610 ;
        RECT 709.285 66.370 713.415 66.670 ;
        RECT 660.325 66.140 692.070 66.160 ;
        RECT 613.575 65.750 619.965 66.040 ;
        RECT 624.845 65.890 692.070 66.140 ;
        RECT 624.845 65.870 660.755 65.890 ;
        RECT 696.290 65.770 702.680 66.060 ;
        RECT 612.990 65.170 623.495 65.505 ;
        RECT 648.465 65.305 659.015 65.640 ;
        RECT 695.705 65.190 706.185 65.525 ;
        RECT 612.340 64.585 615.260 64.885 ;
        RECT 618.805 64.570 622.175 64.870 ;
        RECT 627.055 64.665 628.360 65.045 ;
        RECT 629.060 64.665 632.360 65.045 ;
        RECT 633.060 64.665 636.360 65.045 ;
        RECT 637.060 64.665 638.420 65.045 ;
        RECT 640.395 64.665 641.860 65.045 ;
        RECT 642.560 64.665 645.860 65.045 ;
        RECT 646.560 64.665 649.860 65.045 ;
        RECT 650.560 64.665 651.740 65.045 ;
        RECT 665.675 64.685 666.980 65.065 ;
        RECT 671.680 64.685 674.980 65.065 ;
        RECT 675.680 64.685 677.040 65.065 ;
        RECT 679.015 64.685 680.480 65.065 ;
        RECT 681.180 64.685 684.480 65.065 ;
        RECT 689.180 64.685 690.360 65.065 ;
        RECT 628.520 64.320 628.900 64.355 ;
        RECT 610.555 63.835 610.935 64.215 ;
        RECT 612.960 63.850 614.740 64.140 ;
        RECT 616.215 63.940 617.405 64.225 ;
        RECT 620.335 63.820 621.645 64.140 ;
        RECT 628.255 64.010 631.265 64.320 ;
        RECT 628.520 63.975 628.900 64.010 ;
        RECT 632.520 63.975 633.610 64.355 ;
        RECT 636.520 64.350 636.900 64.355 ;
        RECT 634.040 63.985 636.905 64.350 ;
        RECT 642.020 64.330 642.400 64.355 ;
        RECT 642.005 64.010 644.150 64.330 ;
        RECT 636.520 63.975 636.900 63.985 ;
        RECT 642.020 63.975 642.400 64.010 ;
        RECT 645.065 63.975 646.400 64.355 ;
        RECT 650.020 64.335 650.400 64.355 ;
        RECT 667.140 64.340 667.520 64.375 ;
        RECT 647.555 64.015 650.465 64.335 ;
        RECT 666.875 64.030 669.885 64.340 ;
        RECT 650.020 63.975 650.400 64.015 ;
        RECT 667.140 63.995 667.520 64.030 ;
        RECT 671.140 63.995 672.230 64.375 ;
        RECT 675.140 64.370 675.520 64.375 ;
        RECT 672.660 64.005 675.525 64.370 ;
        RECT 680.640 64.350 681.020 64.375 ;
        RECT 680.625 64.030 682.770 64.350 ;
        RECT 675.140 63.995 675.520 64.005 ;
        RECT 680.640 63.995 681.020 64.030 ;
        RECT 683.685 63.995 685.020 64.375 ;
        RECT 688.640 64.355 689.020 64.375 ;
        RECT 686.175 64.035 689.085 64.355 ;
        RECT 688.640 63.995 689.020 64.035 ;
        RECT 693.270 63.855 693.650 64.235 ;
        RECT 695.675 63.870 697.455 64.160 ;
        RECT 698.930 63.960 700.120 64.245 ;
        RECT 703.050 63.840 704.360 64.160 ;
        RECT 611.690 63.235 612.070 63.615 ;
        RECT 615.435 63.275 615.815 63.655 ;
        RECT 618.145 63.265 618.525 63.645 ;
        RECT 619.555 63.110 622.735 63.430 ;
        RECT 694.405 63.255 694.785 63.635 ;
        RECT 698.150 63.295 698.530 63.675 ;
        RECT 700.860 63.285 701.240 63.665 ;
        RECT 702.270 63.130 705.450 63.450 ;
        RECT 626.870 62.665 628.360 63.045 ;
        RECT 629.060 62.665 630.345 63.045 ;
        RECT 648.375 62.665 649.860 63.045 ;
        RECT 650.560 62.665 651.635 63.045 ;
        RECT 665.490 62.685 666.980 63.065 ;
        RECT 689.180 62.685 690.255 63.065 ;
        RECT 628.520 61.975 629.610 62.355 ;
        RECT 630.565 61.985 632.085 62.345 ;
        RECT 633.005 61.980 645.855 62.315 ;
        RECT 650.020 62.310 650.400 62.355 ;
        RECT 649.285 62.010 650.595 62.310 ;
        RECT 650.020 61.975 650.400 62.010 ;
        RECT 667.140 61.995 668.230 62.375 ;
        RECT 669.185 62.005 670.705 62.365 ;
        RECT 671.625 62.000 684.475 62.335 ;
        RECT 688.640 62.330 689.020 62.375 ;
        RECT 687.905 62.030 689.215 62.330 ;
        RECT 688.640 61.995 689.020 62.030 ;
        RECT 657.700 61.465 690.650 61.500 ;
        RECT 625.375 61.135 690.650 61.465 ;
        RECT 625.375 61.115 658.455 61.135 ;
        RECT 692.445 61.125 696.705 61.480 ;
        RECT 690.650 60.540 696.295 60.545 ;
        RECT 706.910 60.540 707.290 66.370 ;
        RECT 715.790 66.320 720.290 66.630 ;
        RECT 791.990 66.350 796.120 66.650 ;
        RECT 711.750 65.770 718.140 66.060 ;
        RECT 711.165 65.190 727.185 65.525 ;
        RECT 775.835 65.230 781.750 65.565 ;
        RECT 779.105 65.210 781.750 65.230 ;
        RECT 710.515 64.605 713.435 64.905 ;
        RECT 716.980 64.590 720.350 64.890 ;
        RECT 756.430 64.590 759.730 64.970 ;
        RECT 760.430 64.590 763.730 64.970 ;
        RECT 769.930 64.590 773.230 64.970 ;
        RECT 773.930 64.590 777.230 64.970 ;
        RECT 708.730 63.855 709.110 64.235 ;
        RECT 711.135 63.870 712.915 64.160 ;
        RECT 714.390 63.960 715.580 64.245 ;
        RECT 718.510 63.840 719.820 64.160 ;
        RECT 709.865 63.255 710.245 63.635 ;
        RECT 713.610 63.295 713.990 63.675 ;
        RECT 716.320 63.285 716.700 63.665 ;
        RECT 717.730 63.130 720.910 63.450 ;
        RECT 756.430 62.590 757.715 62.970 ;
        RECT 775.745 62.590 777.230 62.970 ;
        RECT 708.010 62.045 712.160 62.315 ;
        RECT 757.935 61.910 759.455 62.270 ;
        RECT 707.660 60.540 711.755 60.545 ;
        RECT 663.995 60.535 696.295 60.540 ;
        RECT 706.540 60.535 711.755 60.540 ;
        RECT 609.485 60.520 613.580 60.525 ;
        RECT 663.995 60.520 721.570 60.535 ;
        RECT 789.615 60.520 789.995 66.350 ;
        RECT 798.495 66.300 802.995 66.610 ;
        RECT 807.450 66.350 811.580 66.650 ;
        RECT 794.455 65.750 800.845 66.040 ;
        RECT 793.870 65.170 804.525 65.505 ;
        RECT 793.220 64.585 796.140 64.885 ;
        RECT 799.685 64.570 803.055 64.870 ;
        RECT 791.435 63.835 791.815 64.215 ;
        RECT 793.840 63.850 795.620 64.140 ;
        RECT 797.095 63.940 798.285 64.225 ;
        RECT 801.215 63.820 802.525 64.140 ;
        RECT 792.570 63.235 792.950 63.615 ;
        RECT 796.315 63.275 796.695 63.655 ;
        RECT 799.025 63.265 799.405 63.645 ;
        RECT 800.435 63.110 803.615 63.430 ;
        RECT 790.365 60.520 794.460 60.525 ;
        RECT 805.075 60.520 805.455 66.350 ;
        RECT 813.955 66.300 818.455 66.610 ;
        RECT 905.625 66.370 909.755 66.670 ;
        RECT 856.665 66.140 888.410 66.160 ;
        RECT 809.915 65.750 816.305 66.040 ;
        RECT 821.185 65.890 888.410 66.140 ;
        RECT 821.185 65.870 857.095 65.890 ;
        RECT 892.630 65.770 899.020 66.060 ;
        RECT 809.330 65.170 819.835 65.505 ;
        RECT 844.805 65.305 855.355 65.640 ;
        RECT 892.045 65.190 902.525 65.525 ;
        RECT 808.680 64.585 811.600 64.885 ;
        RECT 815.145 64.570 818.515 64.870 ;
        RECT 823.395 64.665 824.700 65.045 ;
        RECT 825.400 64.665 828.700 65.045 ;
        RECT 829.400 64.665 832.700 65.045 ;
        RECT 833.400 64.665 834.760 65.045 ;
        RECT 836.735 64.665 838.200 65.045 ;
        RECT 838.900 64.665 842.200 65.045 ;
        RECT 842.900 64.665 846.200 65.045 ;
        RECT 846.900 64.665 848.080 65.045 ;
        RECT 862.015 64.685 863.320 65.065 ;
        RECT 868.020 64.685 871.320 65.065 ;
        RECT 872.020 64.685 873.380 65.065 ;
        RECT 875.355 64.685 876.820 65.065 ;
        RECT 877.520 64.685 880.820 65.065 ;
        RECT 885.520 64.685 886.700 65.065 ;
        RECT 824.860 64.320 825.240 64.355 ;
        RECT 806.895 63.835 807.275 64.215 ;
        RECT 809.300 63.850 811.080 64.140 ;
        RECT 812.555 63.940 813.745 64.225 ;
        RECT 816.675 63.820 817.985 64.140 ;
        RECT 824.595 64.010 827.605 64.320 ;
        RECT 824.860 63.975 825.240 64.010 ;
        RECT 828.860 63.975 829.950 64.355 ;
        RECT 832.860 64.350 833.240 64.355 ;
        RECT 830.380 63.985 833.245 64.350 ;
        RECT 838.360 64.330 838.740 64.355 ;
        RECT 838.345 64.010 840.490 64.330 ;
        RECT 832.860 63.975 833.240 63.985 ;
        RECT 838.360 63.975 838.740 64.010 ;
        RECT 841.405 63.975 842.740 64.355 ;
        RECT 846.360 64.335 846.740 64.355 ;
        RECT 863.480 64.340 863.860 64.375 ;
        RECT 843.895 64.015 846.805 64.335 ;
        RECT 863.215 64.030 866.225 64.340 ;
        RECT 846.360 63.975 846.740 64.015 ;
        RECT 863.480 63.995 863.860 64.030 ;
        RECT 867.480 63.995 868.570 64.375 ;
        RECT 871.480 64.370 871.860 64.375 ;
        RECT 869.000 64.005 871.865 64.370 ;
        RECT 876.980 64.350 877.360 64.375 ;
        RECT 876.965 64.030 879.110 64.350 ;
        RECT 871.480 63.995 871.860 64.005 ;
        RECT 876.980 63.995 877.360 64.030 ;
        RECT 880.025 63.995 881.360 64.375 ;
        RECT 884.980 64.355 885.360 64.375 ;
        RECT 882.515 64.035 885.425 64.355 ;
        RECT 884.980 63.995 885.360 64.035 ;
        RECT 889.610 63.855 889.990 64.235 ;
        RECT 892.015 63.870 893.795 64.160 ;
        RECT 895.270 63.960 896.460 64.245 ;
        RECT 899.390 63.840 900.700 64.160 ;
        RECT 808.030 63.235 808.410 63.615 ;
        RECT 811.775 63.275 812.155 63.655 ;
        RECT 814.485 63.265 814.865 63.645 ;
        RECT 815.895 63.110 819.075 63.430 ;
        RECT 890.745 63.255 891.125 63.635 ;
        RECT 894.490 63.295 894.870 63.675 ;
        RECT 897.200 63.285 897.580 63.665 ;
        RECT 898.610 63.130 901.790 63.450 ;
        RECT 823.210 62.665 824.700 63.045 ;
        RECT 825.400 62.665 826.685 63.045 ;
        RECT 844.715 62.665 846.200 63.045 ;
        RECT 846.900 62.665 847.975 63.045 ;
        RECT 861.830 62.685 863.320 63.065 ;
        RECT 885.520 62.685 886.595 63.065 ;
        RECT 824.860 61.975 825.950 62.355 ;
        RECT 826.905 61.985 828.425 62.345 ;
        RECT 829.345 61.980 842.195 62.315 ;
        RECT 846.360 62.310 846.740 62.355 ;
        RECT 845.625 62.010 846.935 62.310 ;
        RECT 846.360 61.975 846.740 62.010 ;
        RECT 863.480 61.995 864.570 62.375 ;
        RECT 865.525 62.005 867.045 62.365 ;
        RECT 867.965 62.000 880.815 62.335 ;
        RECT 884.980 62.330 885.360 62.375 ;
        RECT 884.245 62.030 885.555 62.330 ;
        RECT 884.980 61.995 885.360 62.030 ;
        RECT 854.040 61.465 886.990 61.500 ;
        RECT 821.715 61.135 886.990 61.465 ;
        RECT 821.715 61.115 854.795 61.135 ;
        RECT 888.785 61.125 893.045 61.480 ;
        RECT 886.990 60.540 892.635 60.545 ;
        RECT 903.250 60.540 903.630 66.370 ;
        RECT 912.130 66.320 916.630 66.630 ;
        RECT 988.330 66.350 992.460 66.650 ;
        RECT 908.090 65.770 914.480 66.060 ;
        RECT 907.505 65.190 923.525 65.525 ;
        RECT 972.220 65.215 978.135 65.550 ;
        RECT 975.490 65.195 978.135 65.215 ;
        RECT 906.855 64.605 909.775 64.905 ;
        RECT 913.320 64.590 916.690 64.890 ;
        RECT 952.815 64.575 956.115 64.955 ;
        RECT 956.815 64.575 960.115 64.955 ;
        RECT 966.315 64.575 969.615 64.955 ;
        RECT 970.315 64.575 973.615 64.955 ;
        RECT 905.070 63.855 905.450 64.235 ;
        RECT 907.475 63.870 909.255 64.160 ;
        RECT 910.730 63.960 911.920 64.245 ;
        RECT 914.850 63.840 916.160 64.160 ;
        RECT 906.205 63.255 906.585 63.635 ;
        RECT 909.950 63.295 910.330 63.675 ;
        RECT 912.660 63.285 913.040 63.665 ;
        RECT 914.070 63.130 917.250 63.450 ;
        RECT 952.815 62.575 954.100 62.955 ;
        RECT 972.130 62.575 973.615 62.955 ;
        RECT 904.350 62.045 908.500 62.315 ;
        RECT 954.320 61.895 955.840 62.255 ;
        RECT 904.000 60.540 908.095 60.545 ;
        RECT 860.335 60.535 892.635 60.540 ;
        RECT 902.880 60.535 908.095 60.540 ;
        RECT 805.825 60.520 809.920 60.525 ;
        RECT 860.335 60.520 917.910 60.535 ;
        RECT 985.955 60.520 986.335 66.350 ;
        RECT 994.835 66.300 999.335 66.610 ;
        RECT 1003.790 66.350 1007.920 66.650 ;
        RECT 990.795 65.750 997.185 66.040 ;
        RECT 990.210 65.170 1000.865 65.505 ;
        RECT 989.560 64.585 992.480 64.885 ;
        RECT 996.025 64.570 999.395 64.870 ;
        RECT 987.775 63.835 988.155 64.215 ;
        RECT 990.180 63.850 991.960 64.140 ;
        RECT 993.435 63.940 994.625 64.225 ;
        RECT 997.555 63.820 998.865 64.140 ;
        RECT 988.910 63.235 989.290 63.615 ;
        RECT 992.655 63.275 993.035 63.655 ;
        RECT 995.365 63.265 995.745 63.645 ;
        RECT 996.775 63.110 999.955 63.430 ;
        RECT 986.705 60.520 990.800 60.525 ;
        RECT 1001.415 60.520 1001.795 66.350 ;
        RECT 1010.295 66.300 1014.795 66.610 ;
        RECT 1101.965 66.370 1106.095 66.670 ;
        RECT 1053.005 66.140 1084.750 66.160 ;
        RECT 1006.255 65.750 1012.645 66.040 ;
        RECT 1017.525 65.890 1084.750 66.140 ;
        RECT 1017.525 65.870 1053.435 65.890 ;
        RECT 1088.970 65.770 1095.360 66.060 ;
        RECT 1005.670 65.170 1016.175 65.505 ;
        RECT 1041.145 65.305 1051.695 65.640 ;
        RECT 1088.385 65.190 1098.865 65.525 ;
        RECT 1005.020 64.585 1007.940 64.885 ;
        RECT 1011.485 64.570 1014.855 64.870 ;
        RECT 1019.735 64.665 1021.040 65.045 ;
        RECT 1021.740 64.665 1025.040 65.045 ;
        RECT 1025.740 64.665 1029.040 65.045 ;
        RECT 1029.740 64.665 1031.100 65.045 ;
        RECT 1033.075 64.665 1034.540 65.045 ;
        RECT 1035.240 64.665 1038.540 65.045 ;
        RECT 1039.240 64.665 1042.540 65.045 ;
        RECT 1043.240 64.665 1044.420 65.045 ;
        RECT 1058.355 64.685 1059.660 65.065 ;
        RECT 1064.360 64.685 1067.660 65.065 ;
        RECT 1068.360 64.685 1069.720 65.065 ;
        RECT 1071.695 64.685 1073.160 65.065 ;
        RECT 1073.860 64.685 1077.160 65.065 ;
        RECT 1081.860 64.685 1083.040 65.065 ;
        RECT 1021.200 64.320 1021.580 64.355 ;
        RECT 1003.235 63.835 1003.615 64.215 ;
        RECT 1005.640 63.850 1007.420 64.140 ;
        RECT 1008.895 63.940 1010.085 64.225 ;
        RECT 1013.015 63.820 1014.325 64.140 ;
        RECT 1020.935 64.010 1023.945 64.320 ;
        RECT 1021.200 63.975 1021.580 64.010 ;
        RECT 1025.200 63.975 1026.290 64.355 ;
        RECT 1029.200 64.350 1029.580 64.355 ;
        RECT 1026.720 63.985 1029.585 64.350 ;
        RECT 1034.700 64.330 1035.080 64.355 ;
        RECT 1034.685 64.010 1036.830 64.330 ;
        RECT 1029.200 63.975 1029.580 63.985 ;
        RECT 1034.700 63.975 1035.080 64.010 ;
        RECT 1037.745 63.975 1039.080 64.355 ;
        RECT 1042.700 64.335 1043.080 64.355 ;
        RECT 1059.820 64.340 1060.200 64.375 ;
        RECT 1040.235 64.015 1043.145 64.335 ;
        RECT 1059.555 64.030 1062.565 64.340 ;
        RECT 1042.700 63.975 1043.080 64.015 ;
        RECT 1059.820 63.995 1060.200 64.030 ;
        RECT 1063.820 63.995 1064.910 64.375 ;
        RECT 1067.820 64.370 1068.200 64.375 ;
        RECT 1065.340 64.005 1068.205 64.370 ;
        RECT 1073.320 64.350 1073.700 64.375 ;
        RECT 1073.305 64.030 1075.450 64.350 ;
        RECT 1067.820 63.995 1068.200 64.005 ;
        RECT 1073.320 63.995 1073.700 64.030 ;
        RECT 1076.365 63.995 1077.700 64.375 ;
        RECT 1081.320 64.355 1081.700 64.375 ;
        RECT 1078.855 64.035 1081.765 64.355 ;
        RECT 1081.320 63.995 1081.700 64.035 ;
        RECT 1085.950 63.855 1086.330 64.235 ;
        RECT 1088.355 63.870 1090.135 64.160 ;
        RECT 1091.610 63.960 1092.800 64.245 ;
        RECT 1095.730 63.840 1097.040 64.160 ;
        RECT 1004.370 63.235 1004.750 63.615 ;
        RECT 1008.115 63.275 1008.495 63.655 ;
        RECT 1010.825 63.265 1011.205 63.645 ;
        RECT 1012.235 63.110 1015.415 63.430 ;
        RECT 1087.085 63.255 1087.465 63.635 ;
        RECT 1090.830 63.295 1091.210 63.675 ;
        RECT 1093.540 63.285 1093.920 63.665 ;
        RECT 1094.950 63.130 1098.130 63.450 ;
        RECT 1019.550 62.665 1021.040 63.045 ;
        RECT 1021.740 62.665 1023.025 63.045 ;
        RECT 1041.055 62.665 1042.540 63.045 ;
        RECT 1043.240 62.665 1044.315 63.045 ;
        RECT 1058.170 62.685 1059.660 63.065 ;
        RECT 1081.860 62.685 1082.935 63.065 ;
        RECT 1021.200 61.975 1022.290 62.355 ;
        RECT 1023.245 61.985 1024.765 62.345 ;
        RECT 1025.685 61.980 1038.535 62.315 ;
        RECT 1042.700 62.310 1043.080 62.355 ;
        RECT 1041.965 62.010 1043.275 62.310 ;
        RECT 1042.700 61.975 1043.080 62.010 ;
        RECT 1059.820 61.995 1060.910 62.375 ;
        RECT 1061.865 62.005 1063.385 62.365 ;
        RECT 1064.305 62.000 1077.155 62.335 ;
        RECT 1081.320 62.330 1081.700 62.375 ;
        RECT 1080.585 62.030 1081.895 62.330 ;
        RECT 1081.320 61.995 1081.700 62.030 ;
        RECT 1050.380 61.465 1083.330 61.500 ;
        RECT 1018.055 61.135 1083.330 61.465 ;
        RECT 1018.055 61.115 1051.135 61.135 ;
        RECT 1085.125 61.125 1089.385 61.480 ;
        RECT 1083.330 60.540 1088.975 60.545 ;
        RECT 1099.590 60.540 1099.970 66.370 ;
        RECT 1108.470 66.320 1112.970 66.630 ;
        RECT 1184.670 66.350 1188.800 66.650 ;
        RECT 1104.430 65.770 1110.820 66.060 ;
        RECT 1103.845 65.190 1119.865 65.525 ;
        RECT 1168.545 65.220 1174.460 65.555 ;
        RECT 1171.815 65.200 1174.460 65.220 ;
        RECT 1103.195 64.605 1106.115 64.905 ;
        RECT 1109.660 64.590 1113.030 64.890 ;
        RECT 1149.140 64.580 1152.440 64.960 ;
        RECT 1153.140 64.580 1156.440 64.960 ;
        RECT 1162.640 64.580 1165.940 64.960 ;
        RECT 1166.640 64.580 1169.940 64.960 ;
        RECT 1101.410 63.855 1101.790 64.235 ;
        RECT 1103.815 63.870 1105.595 64.160 ;
        RECT 1107.070 63.960 1108.260 64.245 ;
        RECT 1111.190 63.840 1112.500 64.160 ;
        RECT 1102.545 63.255 1102.925 63.635 ;
        RECT 1106.290 63.295 1106.670 63.675 ;
        RECT 1109.000 63.285 1109.380 63.665 ;
        RECT 1110.410 63.130 1113.590 63.450 ;
        RECT 1149.140 62.580 1150.425 62.960 ;
        RECT 1168.455 62.580 1169.940 62.960 ;
        RECT 1100.690 62.045 1104.840 62.315 ;
        RECT 1150.645 61.900 1152.165 62.260 ;
        RECT 1100.340 60.540 1104.435 60.545 ;
        RECT 1056.675 60.535 1088.975 60.540 ;
        RECT 1099.220 60.535 1104.435 60.540 ;
        RECT 1002.165 60.520 1006.260 60.525 ;
        RECT 1056.675 60.520 1114.250 60.535 ;
        RECT 1182.295 60.520 1182.675 66.350 ;
        RECT 1191.175 66.300 1195.675 66.610 ;
        RECT 1200.130 66.350 1204.260 66.650 ;
        RECT 1187.135 65.750 1193.525 66.040 ;
        RECT 1186.550 65.170 1197.205 65.505 ;
        RECT 1185.900 64.585 1188.820 64.885 ;
        RECT 1192.365 64.570 1195.735 64.870 ;
        RECT 1184.115 63.835 1184.495 64.215 ;
        RECT 1186.520 63.850 1188.300 64.140 ;
        RECT 1189.775 63.940 1190.965 64.225 ;
        RECT 1193.895 63.820 1195.205 64.140 ;
        RECT 1185.250 63.235 1185.630 63.615 ;
        RECT 1188.995 63.275 1189.375 63.655 ;
        RECT 1191.705 63.265 1192.085 63.645 ;
        RECT 1193.115 63.110 1196.295 63.430 ;
        RECT 1183.045 60.520 1187.140 60.525 ;
        RECT 1197.755 60.520 1198.135 66.350 ;
        RECT 1206.635 66.300 1211.135 66.610 ;
        RECT 1282.845 66.370 1286.975 66.670 ;
        RECT 1289.350 66.320 1293.850 66.630 ;
        RECT 1298.305 66.370 1302.435 66.670 ;
        RECT 1249.345 66.140 1281.090 66.160 ;
        RECT 1202.595 65.750 1208.985 66.040 ;
        RECT 1213.865 65.890 1281.090 66.140 ;
        RECT 1213.865 65.870 1249.775 65.890 ;
        RECT 1285.310 65.770 1291.700 66.060 ;
        RECT 1202.010 65.170 1212.515 65.505 ;
        RECT 1237.485 65.305 1248.035 65.640 ;
        RECT 1276.105 65.325 1280.050 65.660 ;
        RECT 1284.725 65.190 1295.205 65.525 ;
        RECT 1201.360 64.585 1204.280 64.885 ;
        RECT 1207.825 64.570 1211.195 64.870 ;
        RECT 1216.075 64.665 1217.380 65.045 ;
        RECT 1218.080 64.665 1221.380 65.045 ;
        RECT 1222.080 64.665 1225.380 65.045 ;
        RECT 1226.080 64.665 1227.440 65.045 ;
        RECT 1229.415 64.665 1230.880 65.045 ;
        RECT 1231.580 64.665 1234.880 65.045 ;
        RECT 1235.580 64.665 1238.880 65.045 ;
        RECT 1239.580 64.665 1240.760 65.045 ;
        RECT 1254.695 64.685 1256.000 65.065 ;
        RECT 1256.700 64.685 1260.000 65.065 ;
        RECT 1260.700 64.685 1264.000 65.065 ;
        RECT 1264.700 64.685 1266.060 65.065 ;
        RECT 1268.035 64.685 1269.500 65.065 ;
        RECT 1270.200 64.685 1273.500 65.065 ;
        RECT 1274.200 64.685 1277.500 65.065 ;
        RECT 1278.200 64.685 1279.380 65.065 ;
        RECT 1284.075 64.605 1286.995 64.905 ;
        RECT 1290.540 64.590 1293.910 64.890 ;
        RECT 1217.540 64.320 1217.920 64.355 ;
        RECT 1199.575 63.835 1199.955 64.215 ;
        RECT 1201.980 63.850 1203.760 64.140 ;
        RECT 1205.235 63.940 1206.425 64.225 ;
        RECT 1209.355 63.820 1210.665 64.140 ;
        RECT 1217.275 64.010 1220.285 64.320 ;
        RECT 1217.540 63.975 1217.920 64.010 ;
        RECT 1221.540 63.975 1222.630 64.355 ;
        RECT 1225.540 64.350 1225.920 64.355 ;
        RECT 1223.060 63.985 1225.925 64.350 ;
        RECT 1231.040 64.330 1231.420 64.355 ;
        RECT 1231.025 64.010 1233.170 64.330 ;
        RECT 1225.540 63.975 1225.920 63.985 ;
        RECT 1231.040 63.975 1231.420 64.010 ;
        RECT 1234.085 63.975 1235.420 64.355 ;
        RECT 1239.040 64.335 1239.420 64.355 ;
        RECT 1256.160 64.340 1256.540 64.375 ;
        RECT 1236.575 64.015 1239.485 64.335 ;
        RECT 1255.895 64.030 1258.905 64.340 ;
        RECT 1239.040 63.975 1239.420 64.015 ;
        RECT 1256.160 63.995 1256.540 64.030 ;
        RECT 1260.160 63.995 1261.250 64.375 ;
        RECT 1264.160 64.370 1264.540 64.375 ;
        RECT 1261.680 64.005 1264.545 64.370 ;
        RECT 1269.660 64.350 1270.040 64.375 ;
        RECT 1269.645 64.030 1271.790 64.350 ;
        RECT 1264.160 63.995 1264.540 64.005 ;
        RECT 1269.660 63.995 1270.040 64.030 ;
        RECT 1272.705 63.995 1274.040 64.375 ;
        RECT 1277.660 64.355 1278.040 64.375 ;
        RECT 1275.195 64.035 1278.105 64.355 ;
        RECT 1277.660 63.995 1278.040 64.035 ;
        RECT 1282.290 63.855 1282.670 64.235 ;
        RECT 1284.695 63.870 1286.475 64.160 ;
        RECT 1287.950 63.960 1289.140 64.245 ;
        RECT 1292.070 63.840 1293.380 64.160 ;
        RECT 1200.710 63.235 1201.090 63.615 ;
        RECT 1204.455 63.275 1204.835 63.655 ;
        RECT 1207.165 63.265 1207.545 63.645 ;
        RECT 1208.575 63.110 1211.755 63.430 ;
        RECT 1283.425 63.255 1283.805 63.635 ;
        RECT 1287.170 63.295 1287.550 63.675 ;
        RECT 1289.880 63.285 1290.260 63.665 ;
        RECT 1291.290 63.130 1294.470 63.450 ;
        RECT 1215.890 62.665 1217.380 63.045 ;
        RECT 1218.080 62.665 1219.365 63.045 ;
        RECT 1237.395 62.665 1238.880 63.045 ;
        RECT 1239.580 62.665 1240.655 63.045 ;
        RECT 1254.510 62.685 1256.000 63.065 ;
        RECT 1256.700 62.685 1257.985 63.065 ;
        RECT 1276.015 62.685 1277.500 63.065 ;
        RECT 1278.200 62.685 1279.275 63.065 ;
        RECT 1217.540 61.975 1218.630 62.355 ;
        RECT 1219.585 61.985 1221.105 62.345 ;
        RECT 1222.025 61.980 1234.875 62.315 ;
        RECT 1239.040 62.310 1239.420 62.355 ;
        RECT 1238.305 62.010 1239.615 62.310 ;
        RECT 1239.040 61.975 1239.420 62.010 ;
        RECT 1256.160 61.995 1257.250 62.375 ;
        RECT 1258.205 62.005 1259.725 62.365 ;
        RECT 1260.645 62.000 1273.495 62.335 ;
        RECT 1277.660 62.330 1278.040 62.375 ;
        RECT 1276.925 62.030 1278.235 62.330 ;
        RECT 1277.660 61.995 1278.040 62.030 ;
        RECT 1246.720 61.465 1279.670 61.500 ;
        RECT 1214.395 61.135 1279.670 61.465 ;
        RECT 1214.395 61.115 1247.475 61.135 ;
        RECT 1281.465 61.125 1285.725 61.480 ;
        RECT 1279.670 60.540 1285.315 60.545 ;
        RECT 1295.930 60.540 1296.310 66.370 ;
        RECT 1304.810 66.320 1309.310 66.630 ;
        RECT 1300.770 65.770 1307.160 66.060 ;
        RECT 1299.535 64.605 1302.455 64.905 ;
        RECT 1306.000 64.590 1309.370 64.890 ;
        RECT 1297.750 63.855 1298.130 64.235 ;
        RECT 1303.410 63.960 1304.600 64.245 ;
        RECT 1302.630 63.295 1303.010 63.675 ;
        RECT 1306.750 63.130 1309.930 63.450 ;
        RECT 1297.030 62.045 1301.180 62.315 ;
        RECT 1296.680 60.540 1300.775 60.545 ;
        RECT 1253.015 60.535 1285.315 60.540 ;
        RECT 1295.560 60.535 1300.775 60.540 ;
        RECT 1198.505 60.520 1202.600 60.525 ;
        RECT 1253.015 60.520 1310.590 60.535 ;
        RECT 592.905 60.515 598.120 60.520 ;
        RECT 608.365 60.515 613.580 60.520 ;
        RECT 623.825 60.515 721.570 60.520 ;
        RECT 511.285 60.505 515.380 60.510 ;
        RECT 467.620 60.500 499.920 60.505 ;
        RECT 510.165 60.500 515.380 60.505 ;
        RECT 413.110 60.485 417.205 60.490 ;
        RECT 467.620 60.485 525.195 60.500 ;
        RECT 396.530 60.480 401.745 60.485 ;
        RECT 411.990 60.480 417.205 60.485 ;
        RECT 427.450 60.480 525.195 60.485 ;
        RECT 200.130 59.635 271.300 59.655 ;
        RECT 360.060 59.495 386.715 60.395 ;
        RECT 396.530 59.605 525.195 60.480 ;
        RECT 396.530 59.585 467.700 59.605 ;
        RECT 556.380 59.540 583.035 60.440 ;
        RECT 592.905 59.640 721.570 60.515 ;
        RECT 789.245 60.515 794.460 60.520 ;
        RECT 804.705 60.515 809.920 60.520 ;
        RECT 820.165 60.515 917.910 60.520 ;
        RECT 592.905 59.620 664.075 59.640 ;
        RECT 752.745 59.545 779.400 60.445 ;
        RECT 789.245 59.640 917.910 60.515 ;
        RECT 985.585 60.515 990.800 60.520 ;
        RECT 1001.045 60.515 1006.260 60.520 ;
        RECT 1016.505 60.515 1114.250 60.520 ;
        RECT 789.245 59.620 860.415 59.640 ;
        RECT 949.130 59.530 975.785 60.430 ;
        RECT 985.585 59.640 1114.250 60.515 ;
        RECT 1181.925 60.515 1187.140 60.520 ;
        RECT 1197.385 60.515 1202.600 60.520 ;
        RECT 1212.845 60.515 1310.590 60.520 ;
        RECT 985.585 59.620 1056.755 59.640 ;
        RECT 1145.455 59.535 1172.110 60.435 ;
        RECT 1181.925 59.640 1310.590 60.515 ;
        RECT 1181.925 59.620 1253.095 59.640 ;
        RECT -81.535 54.750 -56.100 55.650 ;
        RECT -31.210 54.830 -5.775 55.730 ;
        RECT 3.715 55.610 76.105 55.750 ;
        RECT 3.715 54.850 132.430 55.610 ;
        RECT -79.050 52.570 -77.850 52.950 ;
        RECT -76.095 52.355 -73.820 52.865 ;
        RECT -71.195 52.355 -68.895 52.865 ;
        RECT -66.600 52.355 -64.320 52.865 ;
        RECT -59.525 52.670 -58.290 53.050 ;
        RECT -28.725 52.650 -27.525 53.030 ;
        RECT -25.770 52.435 -23.495 52.945 ;
        RECT -20.870 52.435 -18.570 52.945 ;
        RECT -16.275 52.435 -13.995 52.945 ;
        RECT -9.200 52.750 -7.965 53.130 ;
        RECT -79.050 50.270 -75.790 50.650 ;
        RECT -75.050 50.270 -71.790 50.650 ;
        RECT -65.550 50.270 -62.290 50.650 ;
        RECT -61.550 50.270 -58.290 50.650 ;
        RECT -28.725 50.350 -25.465 50.730 ;
        RECT -24.725 50.350 -21.465 50.730 ;
        RECT -15.225 50.350 -11.965 50.730 ;
        RECT -11.225 50.350 -7.965 50.730 ;
        RECT -78.385 48.685 -56.100 48.695 ;
        RECT -78.385 48.355 -54.560 48.685 ;
        RECT -28.060 48.435 -1.765 48.775 ;
        RECT -56.320 48.335 -54.560 48.355 ;
        RECT 4.085 47.690 4.465 54.850 ;
        RECT 5.915 50.635 9.290 51.035 ;
        RECT 9.660 50.395 10.040 50.775 ;
        RECT 12.375 50.435 12.755 50.815 ;
        RECT 16.560 50.385 16.940 50.765 ;
        RECT 6.985 49.970 8.725 50.260 ;
        RECT 10.775 49.920 11.975 50.210 ;
        RECT 13.485 49.890 16.095 50.315 ;
        RECT 17.695 49.985 18.075 50.365 ;
        RECT 5.230 49.210 18.795 49.525 ;
        RECT 5.225 48.465 18.785 48.765 ;
        RECT 5.245 47.750 11.970 48.050 ;
        RECT 15.670 47.450 18.775 47.725 ;
        RECT 19.545 47.690 19.925 54.850 ;
        RECT 76.075 54.710 132.430 54.850 ;
        RECT 164.960 54.840 190.395 55.740 ;
        RECT 200.080 55.610 272.470 55.750 ;
        RECT 200.080 54.850 328.795 55.610 ;
        RECT 36.185 53.725 73.735 53.865 ;
        RECT 36.185 53.580 101.835 53.725 ;
        RECT 73.060 53.440 101.835 53.580 ;
        RECT 103.505 53.420 110.210 53.720 ;
        RECT 37.695 52.670 39.150 53.050 ;
        RECT 39.890 52.670 41.090 53.050 ;
        RECT 42.845 52.455 45.120 52.965 ;
        RECT 47.745 52.455 50.045 52.965 ;
        RECT 52.340 52.455 54.620 52.965 ;
        RECT 59.415 52.770 60.650 53.150 ;
        RECT 61.390 52.770 62.670 53.150 ;
        RECT 76.365 52.530 77.820 52.910 ;
        RECT 60.830 52.415 61.210 52.450 ;
        RECT 39.330 52.310 39.710 52.350 ;
        RECT 39.260 52.005 42.095 52.310 ;
        RECT 58.075 52.105 61.210 52.415 ;
        RECT 81.515 52.315 83.790 52.825 ;
        RECT 86.415 52.315 88.715 52.825 ;
        RECT 91.010 52.315 93.290 52.825 ;
        RECT 100.060 52.630 101.340 53.010 ;
        RECT 99.500 52.275 99.880 52.310 ;
        RECT 78.000 52.170 78.380 52.210 ;
        RECT 60.830 52.070 61.210 52.105 ;
        RECT 39.330 51.970 39.710 52.005 ;
        RECT 77.930 51.865 80.765 52.170 ;
        RECT 96.745 51.965 99.880 52.275 ;
        RECT 99.500 51.930 99.880 51.965 ;
        RECT 78.000 51.830 78.380 51.865 ;
        RECT 21.375 50.595 24.780 51.035 ;
        RECT 25.120 50.395 25.500 50.775 ;
        RECT 27.835 50.435 28.215 50.815 ;
        RECT 32.020 50.385 32.400 50.765 ;
        RECT 37.855 50.370 39.150 50.750 ;
        RECT 39.890 50.370 43.150 50.750 ;
        RECT 43.890 50.370 47.150 50.750 ;
        RECT 47.890 50.370 49.075 50.750 ;
        RECT 51.340 50.370 52.650 50.750 ;
        RECT 53.390 50.370 56.650 50.750 ;
        RECT 57.390 50.370 60.650 50.750 ;
        RECT 61.390 50.370 62.405 50.750 ;
        RECT 22.445 49.970 24.185 50.260 ;
        RECT 26.235 49.920 27.435 50.210 ;
        RECT 28.945 49.890 31.540 50.265 ;
        RECT 33.155 49.985 33.535 50.365 ;
        RECT 76.525 50.230 77.820 50.610 ;
        RECT 82.560 50.230 85.820 50.610 ;
        RECT 86.560 50.230 87.745 50.610 ;
        RECT 90.010 50.230 91.320 50.610 ;
        RECT 92.060 50.230 95.320 50.610 ;
        RECT 100.060 50.230 101.075 50.610 ;
        RECT 104.140 50.475 107.555 50.895 ;
        RECT 107.885 50.255 108.265 50.635 ;
        RECT 110.600 50.295 110.980 50.675 ;
        RECT 114.785 50.245 115.165 50.625 ;
        RECT 39.330 49.670 39.710 50.050 ;
        RECT 43.330 49.670 43.710 50.050 ;
        RECT 47.330 50.005 47.710 50.050 ;
        RECT 52.830 50.005 53.210 50.050 ;
        RECT 47.280 49.690 53.215 50.005 ;
        RECT 47.330 49.670 47.710 49.690 ;
        RECT 52.830 49.670 53.210 49.690 ;
        RECT 56.830 49.670 57.210 50.050 ;
        RECT 60.830 49.670 61.210 50.050 ;
        RECT 78.000 49.530 78.380 49.910 ;
        RECT 82.000 49.530 82.380 49.910 ;
        RECT 86.000 49.865 86.380 49.910 ;
        RECT 91.500 49.865 91.880 49.910 ;
        RECT 85.950 49.550 91.885 49.865 ;
        RECT 86.000 49.530 86.380 49.550 ;
        RECT 91.500 49.530 91.880 49.550 ;
        RECT 95.500 49.530 95.880 49.910 ;
        RECT 99.500 49.530 99.880 49.910 ;
        RECT 105.210 49.830 106.950 50.120 ;
        RECT 109.000 49.780 110.200 50.070 ;
        RECT 111.710 49.740 114.340 50.195 ;
        RECT 115.920 49.845 116.300 50.225 ;
        RECT 20.685 49.210 34.510 49.510 ;
        RECT 36.185 49.045 52.195 49.420 ;
        RECT 70.090 48.905 90.865 49.280 ;
        RECT 20.690 48.465 39.110 48.765 ;
        RECT 40.555 48.455 67.865 48.795 ;
        RECT 20.170 47.750 27.430 48.050 ;
        RECT 5.225 47.130 9.350 47.400 ;
        RECT 20.725 47.215 24.810 47.485 ;
        RECT 31.130 47.450 34.880 47.725 ;
        RECT 36.185 47.690 62.415 48.080 ;
        RECT 69.120 47.550 101.085 47.940 ;
        RECT 36.185 47.325 54.855 47.335 ;
        RECT 36.185 47.195 66.205 47.325 ;
        RECT 113.895 47.310 117.025 47.585 ;
        RECT 117.770 47.550 118.150 54.710 ;
        RECT 167.445 52.660 168.645 53.040 ;
        RECT 119.010 52.250 125.750 52.550 ;
        RECT 170.400 52.445 172.675 52.955 ;
        RECT 175.300 52.445 177.600 52.955 ;
        RECT 179.895 52.445 182.175 52.955 ;
        RECT 186.970 52.760 188.205 53.140 ;
        RECT 119.600 50.455 123.055 50.895 ;
        RECT 123.345 50.255 123.725 50.635 ;
        RECT 126.060 50.295 126.440 50.675 ;
        RECT 130.245 50.245 130.625 50.625 ;
        RECT 167.445 50.360 170.705 50.740 ;
        RECT 171.445 50.360 174.705 50.740 ;
        RECT 180.945 50.360 184.205 50.740 ;
        RECT 184.945 50.360 188.205 50.740 ;
        RECT 120.670 49.830 122.410 50.120 ;
        RECT 124.460 49.780 125.660 50.070 ;
        RECT 127.170 49.750 129.795 50.160 ;
        RECT 131.380 49.845 131.760 50.225 ;
        RECT 118.415 49.070 134.335 49.370 ;
        RECT 118.950 48.325 135.895 48.625 ;
        RECT 168.110 48.445 194.405 48.785 ;
        RECT 200.450 47.690 200.830 54.850 ;
        RECT 202.280 50.635 205.655 51.035 ;
        RECT 206.025 50.395 206.405 50.775 ;
        RECT 208.740 50.435 209.120 50.815 ;
        RECT 212.925 50.385 213.305 50.765 ;
        RECT 203.350 49.970 205.090 50.260 ;
        RECT 207.140 49.920 208.340 50.210 ;
        RECT 209.850 49.890 212.460 50.315 ;
        RECT 214.060 49.985 214.440 50.365 ;
        RECT 201.595 49.210 215.160 49.525 ;
        RECT 201.590 48.465 215.150 48.765 ;
        RECT 201.610 47.750 208.335 48.050 ;
        RECT 129.355 47.310 137.055 47.585 ;
        RECT 212.035 47.450 215.140 47.725 ;
        RECT 215.910 47.690 216.290 54.850 ;
        RECT 272.440 54.710 328.795 54.850 ;
        RECT 361.350 54.800 386.785 55.700 ;
        RECT 396.480 55.560 468.870 55.700 ;
        RECT 396.480 54.800 525.195 55.560 ;
        RECT 557.670 54.845 583.105 55.745 ;
        RECT 592.855 55.595 665.245 55.735 ;
        RECT 592.855 54.835 721.570 55.595 ;
        RECT 754.035 54.850 779.470 55.750 ;
        RECT 789.195 55.595 861.585 55.735 ;
        RECT 789.195 54.835 917.910 55.595 ;
        RECT 950.420 54.835 975.855 55.735 ;
        RECT 985.535 55.595 1057.925 55.735 ;
        RECT 985.535 54.835 1114.250 55.595 ;
        RECT 1146.745 54.840 1172.180 55.740 ;
        RECT 1181.875 55.595 1254.265 55.735 ;
        RECT 1181.875 54.835 1310.590 55.595 ;
        RECT 232.550 53.725 270.100 53.865 ;
        RECT 232.550 53.580 298.200 53.725 ;
        RECT 269.425 53.440 298.200 53.580 ;
        RECT 299.870 53.420 306.575 53.720 ;
        RECT 234.060 52.670 235.515 53.050 ;
        RECT 236.255 52.670 237.455 53.050 ;
        RECT 239.210 52.455 241.485 52.965 ;
        RECT 244.110 52.455 246.410 52.965 ;
        RECT 248.705 52.455 250.985 52.965 ;
        RECT 255.780 52.770 257.015 53.150 ;
        RECT 257.755 52.770 259.035 53.150 ;
        RECT 272.730 52.530 274.185 52.910 ;
        RECT 257.195 52.415 257.575 52.450 ;
        RECT 235.695 52.310 236.075 52.350 ;
        RECT 235.625 52.005 238.460 52.310 ;
        RECT 254.440 52.105 257.575 52.415 ;
        RECT 277.880 52.315 280.155 52.825 ;
        RECT 282.780 52.315 285.080 52.825 ;
        RECT 287.375 52.315 289.655 52.825 ;
        RECT 296.425 52.630 297.705 53.010 ;
        RECT 295.865 52.275 296.245 52.310 ;
        RECT 274.365 52.170 274.745 52.210 ;
        RECT 257.195 52.070 257.575 52.105 ;
        RECT 235.695 51.970 236.075 52.005 ;
        RECT 274.295 51.865 277.130 52.170 ;
        RECT 293.110 51.965 296.245 52.275 ;
        RECT 295.865 51.930 296.245 51.965 ;
        RECT 274.365 51.830 274.745 51.865 ;
        RECT 217.740 50.595 221.145 51.035 ;
        RECT 221.485 50.395 221.865 50.775 ;
        RECT 224.200 50.435 224.580 50.815 ;
        RECT 228.385 50.385 228.765 50.765 ;
        RECT 234.220 50.370 235.515 50.750 ;
        RECT 236.255 50.370 239.515 50.750 ;
        RECT 240.255 50.370 243.515 50.750 ;
        RECT 244.255 50.370 245.440 50.750 ;
        RECT 247.705 50.370 249.015 50.750 ;
        RECT 249.755 50.370 253.015 50.750 ;
        RECT 253.755 50.370 257.015 50.750 ;
        RECT 257.755 50.370 258.770 50.750 ;
        RECT 218.810 49.970 220.550 50.260 ;
        RECT 222.600 49.920 223.800 50.210 ;
        RECT 225.310 49.890 227.905 50.265 ;
        RECT 229.520 49.985 229.900 50.365 ;
        RECT 272.890 50.230 274.185 50.610 ;
        RECT 278.925 50.230 282.185 50.610 ;
        RECT 282.925 50.230 284.110 50.610 ;
        RECT 286.375 50.230 287.685 50.610 ;
        RECT 288.425 50.230 291.685 50.610 ;
        RECT 296.425 50.230 297.440 50.610 ;
        RECT 300.505 50.475 303.920 50.895 ;
        RECT 304.250 50.255 304.630 50.635 ;
        RECT 306.965 50.295 307.345 50.675 ;
        RECT 311.150 50.245 311.530 50.625 ;
        RECT 235.695 49.670 236.075 50.050 ;
        RECT 239.695 49.670 240.075 50.050 ;
        RECT 243.695 50.005 244.075 50.050 ;
        RECT 249.195 50.005 249.575 50.050 ;
        RECT 243.645 49.690 249.580 50.005 ;
        RECT 243.695 49.670 244.075 49.690 ;
        RECT 249.195 49.670 249.575 49.690 ;
        RECT 253.195 49.670 253.575 50.050 ;
        RECT 257.195 49.670 257.575 50.050 ;
        RECT 274.365 49.530 274.745 49.910 ;
        RECT 278.365 49.530 278.745 49.910 ;
        RECT 282.365 49.865 282.745 49.910 ;
        RECT 287.865 49.865 288.245 49.910 ;
        RECT 282.315 49.550 288.250 49.865 ;
        RECT 282.365 49.530 282.745 49.550 ;
        RECT 287.865 49.530 288.245 49.550 ;
        RECT 291.865 49.530 292.245 49.910 ;
        RECT 295.865 49.530 296.245 49.910 ;
        RECT 301.575 49.830 303.315 50.120 ;
        RECT 305.365 49.780 306.565 50.070 ;
        RECT 308.075 49.740 310.705 50.195 ;
        RECT 312.285 49.845 312.665 50.225 ;
        RECT 217.050 49.210 230.875 49.510 ;
        RECT 232.550 49.045 248.560 49.420 ;
        RECT 266.455 48.905 287.230 49.280 ;
        RECT 217.055 48.465 235.475 48.765 ;
        RECT 236.920 48.455 264.230 48.795 ;
        RECT 216.535 47.750 223.795 48.050 ;
        RECT 36.185 47.185 93.525 47.195 ;
        RECT 36.185 47.015 102.530 47.185 ;
        RECT 201.590 47.130 205.715 47.400 ;
        RECT 217.090 47.215 221.175 47.485 ;
        RECT 227.495 47.450 231.245 47.725 ;
        RECT 232.550 47.690 258.780 48.080 ;
        RECT 265.485 47.550 297.450 47.940 ;
        RECT 232.550 47.325 251.220 47.335 ;
        RECT 232.550 47.195 262.570 47.325 ;
        RECT 310.260 47.310 313.390 47.585 ;
        RECT 314.135 47.550 314.515 54.710 ;
        RECT 363.835 52.620 365.035 53.000 ;
        RECT 315.375 52.250 322.115 52.550 ;
        RECT 366.790 52.405 369.065 52.915 ;
        RECT 371.690 52.405 373.990 52.915 ;
        RECT 376.285 52.405 378.565 52.915 ;
        RECT 383.360 52.720 384.595 53.100 ;
        RECT 315.965 50.455 319.420 50.895 ;
        RECT 319.710 50.255 320.090 50.635 ;
        RECT 322.425 50.295 322.805 50.675 ;
        RECT 326.610 50.245 326.990 50.625 ;
        RECT 363.835 50.320 367.095 50.700 ;
        RECT 367.835 50.320 371.095 50.700 ;
        RECT 377.335 50.320 380.595 50.700 ;
        RECT 381.335 50.320 384.595 50.700 ;
        RECT 317.035 49.830 318.775 50.120 ;
        RECT 320.825 49.780 322.025 50.070 ;
        RECT 323.535 49.750 326.160 50.160 ;
        RECT 327.745 49.845 328.125 50.225 ;
        RECT 314.780 49.070 330.700 49.370 ;
        RECT 315.315 48.325 332.260 48.625 ;
        RECT 364.500 48.405 390.795 48.745 ;
        RECT 396.850 47.640 397.230 54.800 ;
        RECT 398.680 50.585 402.055 50.985 ;
        RECT 402.425 50.345 402.805 50.725 ;
        RECT 405.140 50.385 405.520 50.765 ;
        RECT 409.325 50.335 409.705 50.715 ;
        RECT 399.750 49.920 401.490 50.210 ;
        RECT 403.540 49.870 404.740 50.160 ;
        RECT 406.250 49.840 408.860 50.265 ;
        RECT 410.460 49.935 410.840 50.315 ;
        RECT 397.995 49.160 411.560 49.475 ;
        RECT 397.990 48.415 411.550 48.715 ;
        RECT 398.010 47.700 404.735 48.000 ;
        RECT 325.720 47.310 333.420 47.585 ;
        RECT 408.435 47.400 411.540 47.675 ;
        RECT 412.310 47.640 412.690 54.800 ;
        RECT 468.840 54.660 525.195 54.800 ;
        RECT 428.950 53.675 466.500 53.815 ;
        RECT 428.950 53.530 494.600 53.675 ;
        RECT 465.825 53.390 494.600 53.530 ;
        RECT 496.270 53.370 502.975 53.670 ;
        RECT 430.460 52.620 431.915 53.000 ;
        RECT 432.655 52.620 433.855 53.000 ;
        RECT 435.610 52.405 437.885 52.915 ;
        RECT 440.510 52.405 442.810 52.915 ;
        RECT 445.105 52.405 447.385 52.915 ;
        RECT 452.180 52.720 453.415 53.100 ;
        RECT 454.155 52.720 455.435 53.100 ;
        RECT 469.130 52.480 470.585 52.860 ;
        RECT 453.595 52.365 453.975 52.400 ;
        RECT 432.095 52.260 432.475 52.300 ;
        RECT 432.025 51.955 434.860 52.260 ;
        RECT 450.840 52.055 453.975 52.365 ;
        RECT 474.280 52.265 476.555 52.775 ;
        RECT 479.180 52.265 481.480 52.775 ;
        RECT 483.775 52.265 486.055 52.775 ;
        RECT 492.825 52.580 494.105 52.960 ;
        RECT 492.265 52.225 492.645 52.260 ;
        RECT 470.765 52.120 471.145 52.160 ;
        RECT 453.595 52.020 453.975 52.055 ;
        RECT 432.095 51.920 432.475 51.955 ;
        RECT 470.695 51.815 473.530 52.120 ;
        RECT 489.510 51.915 492.645 52.225 ;
        RECT 492.265 51.880 492.645 51.915 ;
        RECT 470.765 51.780 471.145 51.815 ;
        RECT 414.140 50.545 417.545 50.985 ;
        RECT 417.885 50.345 418.265 50.725 ;
        RECT 420.600 50.385 420.980 50.765 ;
        RECT 424.785 50.335 425.165 50.715 ;
        RECT 430.620 50.320 431.915 50.700 ;
        RECT 432.655 50.320 435.915 50.700 ;
        RECT 436.655 50.320 439.915 50.700 ;
        RECT 440.655 50.320 441.840 50.700 ;
        RECT 444.105 50.320 445.415 50.700 ;
        RECT 446.155 50.320 449.415 50.700 ;
        RECT 450.155 50.320 453.415 50.700 ;
        RECT 454.155 50.320 455.170 50.700 ;
        RECT 415.210 49.920 416.950 50.210 ;
        RECT 419.000 49.870 420.200 50.160 ;
        RECT 421.710 49.840 424.305 50.215 ;
        RECT 425.920 49.935 426.300 50.315 ;
        RECT 469.290 50.180 470.585 50.560 ;
        RECT 475.325 50.180 478.585 50.560 ;
        RECT 479.325 50.180 480.510 50.560 ;
        RECT 482.775 50.180 484.085 50.560 ;
        RECT 484.825 50.180 488.085 50.560 ;
        RECT 492.825 50.180 493.840 50.560 ;
        RECT 496.905 50.425 500.320 50.845 ;
        RECT 500.650 50.205 501.030 50.585 ;
        RECT 503.365 50.245 503.745 50.625 ;
        RECT 507.550 50.195 507.930 50.575 ;
        RECT 432.095 49.620 432.475 50.000 ;
        RECT 436.095 49.620 436.475 50.000 ;
        RECT 440.095 49.955 440.475 50.000 ;
        RECT 445.595 49.955 445.975 50.000 ;
        RECT 440.045 49.640 445.980 49.955 ;
        RECT 440.095 49.620 440.475 49.640 ;
        RECT 445.595 49.620 445.975 49.640 ;
        RECT 449.595 49.620 449.975 50.000 ;
        RECT 453.595 49.620 453.975 50.000 ;
        RECT 470.765 49.480 471.145 49.860 ;
        RECT 474.765 49.480 475.145 49.860 ;
        RECT 478.765 49.815 479.145 49.860 ;
        RECT 484.265 49.815 484.645 49.860 ;
        RECT 478.715 49.500 484.650 49.815 ;
        RECT 478.765 49.480 479.145 49.500 ;
        RECT 484.265 49.480 484.645 49.500 ;
        RECT 488.265 49.480 488.645 49.860 ;
        RECT 492.265 49.480 492.645 49.860 ;
        RECT 497.975 49.780 499.715 50.070 ;
        RECT 501.765 49.730 502.965 50.020 ;
        RECT 504.475 49.690 507.105 50.145 ;
        RECT 508.685 49.795 509.065 50.175 ;
        RECT 413.450 49.160 427.275 49.460 ;
        RECT 428.950 48.995 444.960 49.370 ;
        RECT 462.855 48.855 483.630 49.230 ;
        RECT 413.455 48.415 431.875 48.715 ;
        RECT 433.320 48.405 460.630 48.745 ;
        RECT 412.935 47.700 420.195 48.000 ;
        RECT 232.550 47.185 289.890 47.195 ;
        RECT 232.550 47.015 298.895 47.185 ;
        RECT 397.990 47.080 402.115 47.350 ;
        RECT 413.490 47.165 417.575 47.435 ;
        RECT 423.895 47.400 427.645 47.675 ;
        RECT 428.950 47.640 455.180 48.030 ;
        RECT 461.885 47.500 493.850 47.890 ;
        RECT 428.950 47.275 447.620 47.285 ;
        RECT 428.950 47.145 458.970 47.275 ;
        RECT 506.660 47.260 509.790 47.535 ;
        RECT 510.535 47.500 510.915 54.660 ;
        RECT 560.155 52.665 561.355 53.045 ;
        RECT 511.775 52.200 518.515 52.500 ;
        RECT 563.110 52.450 565.385 52.960 ;
        RECT 568.010 52.450 570.310 52.960 ;
        RECT 572.605 52.450 574.885 52.960 ;
        RECT 579.680 52.765 580.915 53.145 ;
        RECT 512.365 50.405 515.820 50.845 ;
        RECT 516.110 50.205 516.490 50.585 ;
        RECT 518.825 50.245 519.205 50.625 ;
        RECT 523.010 50.195 523.390 50.575 ;
        RECT 560.155 50.365 563.415 50.745 ;
        RECT 564.155 50.365 567.415 50.745 ;
        RECT 573.655 50.365 576.915 50.745 ;
        RECT 577.655 50.365 580.915 50.745 ;
        RECT 513.435 49.780 515.175 50.070 ;
        RECT 517.225 49.730 518.425 50.020 ;
        RECT 519.935 49.700 522.560 50.110 ;
        RECT 524.145 49.795 524.525 50.175 ;
        RECT 511.180 49.020 527.100 49.320 ;
        RECT 511.715 48.275 528.660 48.575 ;
        RECT 560.820 48.450 587.115 48.790 ;
        RECT 593.225 47.675 593.605 54.835 ;
        RECT 595.055 50.620 598.430 51.020 ;
        RECT 598.800 50.380 599.180 50.760 ;
        RECT 601.515 50.420 601.895 50.800 ;
        RECT 605.700 50.370 606.080 50.750 ;
        RECT 596.125 49.955 597.865 50.245 ;
        RECT 599.915 49.905 601.115 50.195 ;
        RECT 602.625 49.875 605.235 50.300 ;
        RECT 606.835 49.970 607.215 50.350 ;
        RECT 594.370 49.195 607.935 49.510 ;
        RECT 594.365 48.450 607.925 48.750 ;
        RECT 594.385 47.735 601.110 48.035 ;
        RECT 522.120 47.260 529.820 47.535 ;
        RECT 604.810 47.435 607.915 47.710 ;
        RECT 608.685 47.675 609.065 54.835 ;
        RECT 665.215 54.695 721.570 54.835 ;
        RECT 625.325 53.710 662.875 53.850 ;
        RECT 625.325 53.565 690.975 53.710 ;
        RECT 662.200 53.425 690.975 53.565 ;
        RECT 692.645 53.405 699.350 53.705 ;
        RECT 626.835 52.655 628.290 53.035 ;
        RECT 629.030 52.655 630.230 53.035 ;
        RECT 631.985 52.440 634.260 52.950 ;
        RECT 636.885 52.440 639.185 52.950 ;
        RECT 641.480 52.440 643.760 52.950 ;
        RECT 648.555 52.755 649.790 53.135 ;
        RECT 650.530 52.755 651.810 53.135 ;
        RECT 665.505 52.515 666.960 52.895 ;
        RECT 649.970 52.400 650.350 52.435 ;
        RECT 628.470 52.295 628.850 52.335 ;
        RECT 628.400 51.990 631.235 52.295 ;
        RECT 647.215 52.090 650.350 52.400 ;
        RECT 670.655 52.300 672.930 52.810 ;
        RECT 675.555 52.300 677.855 52.810 ;
        RECT 680.150 52.300 682.430 52.810 ;
        RECT 689.200 52.615 690.480 52.995 ;
        RECT 688.640 52.260 689.020 52.295 ;
        RECT 667.140 52.155 667.520 52.195 ;
        RECT 649.970 52.055 650.350 52.090 ;
        RECT 628.470 51.955 628.850 51.990 ;
        RECT 667.070 51.850 669.905 52.155 ;
        RECT 685.885 51.950 689.020 52.260 ;
        RECT 688.640 51.915 689.020 51.950 ;
        RECT 667.140 51.815 667.520 51.850 ;
        RECT 610.515 50.580 613.920 51.020 ;
        RECT 614.260 50.380 614.640 50.760 ;
        RECT 616.975 50.420 617.355 50.800 ;
        RECT 621.160 50.370 621.540 50.750 ;
        RECT 626.995 50.355 628.290 50.735 ;
        RECT 629.030 50.355 632.290 50.735 ;
        RECT 633.030 50.355 636.290 50.735 ;
        RECT 637.030 50.355 638.215 50.735 ;
        RECT 640.480 50.355 641.790 50.735 ;
        RECT 642.530 50.355 645.790 50.735 ;
        RECT 646.530 50.355 649.790 50.735 ;
        RECT 650.530 50.355 651.545 50.735 ;
        RECT 611.585 49.955 613.325 50.245 ;
        RECT 615.375 49.905 616.575 50.195 ;
        RECT 618.085 49.875 620.680 50.250 ;
        RECT 622.295 49.970 622.675 50.350 ;
        RECT 665.665 50.215 666.960 50.595 ;
        RECT 671.700 50.215 674.960 50.595 ;
        RECT 675.700 50.215 676.885 50.595 ;
        RECT 679.150 50.215 680.460 50.595 ;
        RECT 681.200 50.215 684.460 50.595 ;
        RECT 689.200 50.215 690.215 50.595 ;
        RECT 693.280 50.460 696.695 50.880 ;
        RECT 697.025 50.240 697.405 50.620 ;
        RECT 699.740 50.280 700.120 50.660 ;
        RECT 703.925 50.230 704.305 50.610 ;
        RECT 628.470 49.655 628.850 50.035 ;
        RECT 632.470 49.655 632.850 50.035 ;
        RECT 636.470 49.990 636.850 50.035 ;
        RECT 641.970 49.990 642.350 50.035 ;
        RECT 636.420 49.675 642.355 49.990 ;
        RECT 636.470 49.655 636.850 49.675 ;
        RECT 641.970 49.655 642.350 49.675 ;
        RECT 645.970 49.655 646.350 50.035 ;
        RECT 649.970 49.655 650.350 50.035 ;
        RECT 667.140 49.515 667.520 49.895 ;
        RECT 671.140 49.515 671.520 49.895 ;
        RECT 675.140 49.850 675.520 49.895 ;
        RECT 680.640 49.850 681.020 49.895 ;
        RECT 675.090 49.535 681.025 49.850 ;
        RECT 675.140 49.515 675.520 49.535 ;
        RECT 680.640 49.515 681.020 49.535 ;
        RECT 684.640 49.515 685.020 49.895 ;
        RECT 688.640 49.515 689.020 49.895 ;
        RECT 694.350 49.815 696.090 50.105 ;
        RECT 698.140 49.765 699.340 50.055 ;
        RECT 700.850 49.725 703.480 50.180 ;
        RECT 705.060 49.830 705.440 50.210 ;
        RECT 609.825 49.195 623.650 49.495 ;
        RECT 625.325 49.030 641.335 49.405 ;
        RECT 659.230 48.890 680.005 49.265 ;
        RECT 609.830 48.450 628.250 48.750 ;
        RECT 629.695 48.440 657.005 48.780 ;
        RECT 609.310 47.735 616.570 48.035 ;
        RECT 428.950 47.135 486.290 47.145 ;
        RECT 65.965 46.875 102.530 47.015 ;
        RECT 262.330 46.875 298.895 47.015 ;
        RECT 428.950 46.965 495.295 47.135 ;
        RECT 594.365 47.115 598.490 47.385 ;
        RECT 609.865 47.200 613.950 47.470 ;
        RECT 620.270 47.435 624.020 47.710 ;
        RECT 625.325 47.675 651.555 48.065 ;
        RECT 658.260 47.535 690.225 47.925 ;
        RECT 625.325 47.310 643.995 47.320 ;
        RECT 625.325 47.180 655.345 47.310 ;
        RECT 703.035 47.295 706.165 47.570 ;
        RECT 706.910 47.535 707.290 54.695 ;
        RECT 756.520 52.670 757.720 53.050 ;
        RECT 708.150 52.235 714.890 52.535 ;
        RECT 759.475 52.455 761.750 52.965 ;
        RECT 764.375 52.455 766.675 52.965 ;
        RECT 768.970 52.455 771.250 52.965 ;
        RECT 776.045 52.770 777.280 53.150 ;
        RECT 708.740 50.440 712.195 50.880 ;
        RECT 712.485 50.240 712.865 50.620 ;
        RECT 715.200 50.280 715.580 50.660 ;
        RECT 719.385 50.230 719.765 50.610 ;
        RECT 756.520 50.370 759.780 50.750 ;
        RECT 760.520 50.370 763.780 50.750 ;
        RECT 770.020 50.370 773.280 50.750 ;
        RECT 774.020 50.370 777.280 50.750 ;
        RECT 709.810 49.815 711.550 50.105 ;
        RECT 713.600 49.765 714.800 50.055 ;
        RECT 716.310 49.735 718.935 50.145 ;
        RECT 720.520 49.830 720.900 50.210 ;
        RECT 707.555 49.055 723.475 49.355 ;
        RECT 708.090 48.310 725.035 48.610 ;
        RECT 757.185 48.455 783.480 48.795 ;
        RECT 789.565 47.675 789.945 54.835 ;
        RECT 791.395 50.620 794.770 51.020 ;
        RECT 795.140 50.380 795.520 50.760 ;
        RECT 797.855 50.420 798.235 50.800 ;
        RECT 802.040 50.370 802.420 50.750 ;
        RECT 792.465 49.955 794.205 50.245 ;
        RECT 796.255 49.905 797.455 50.195 ;
        RECT 798.965 49.875 801.575 50.300 ;
        RECT 803.175 49.970 803.555 50.350 ;
        RECT 790.710 49.195 804.275 49.510 ;
        RECT 790.705 48.450 804.265 48.750 ;
        RECT 790.725 47.735 797.450 48.035 ;
        RECT 718.495 47.295 726.195 47.570 ;
        RECT 801.150 47.435 804.255 47.710 ;
        RECT 805.025 47.675 805.405 54.835 ;
        RECT 861.555 54.695 917.910 54.835 ;
        RECT 821.665 53.710 859.215 53.850 ;
        RECT 821.665 53.565 887.315 53.710 ;
        RECT 858.540 53.425 887.315 53.565 ;
        RECT 888.985 53.405 895.690 53.705 ;
        RECT 823.175 52.655 824.630 53.035 ;
        RECT 825.370 52.655 826.570 53.035 ;
        RECT 828.325 52.440 830.600 52.950 ;
        RECT 833.225 52.440 835.525 52.950 ;
        RECT 837.820 52.440 840.100 52.950 ;
        RECT 844.895 52.755 846.130 53.135 ;
        RECT 846.870 52.755 848.150 53.135 ;
        RECT 861.845 52.515 863.300 52.895 ;
        RECT 846.310 52.400 846.690 52.435 ;
        RECT 824.810 52.295 825.190 52.335 ;
        RECT 824.740 51.990 827.575 52.295 ;
        RECT 843.555 52.090 846.690 52.400 ;
        RECT 866.995 52.300 869.270 52.810 ;
        RECT 871.895 52.300 874.195 52.810 ;
        RECT 876.490 52.300 878.770 52.810 ;
        RECT 885.540 52.615 886.820 52.995 ;
        RECT 884.980 52.260 885.360 52.295 ;
        RECT 863.480 52.155 863.860 52.195 ;
        RECT 846.310 52.055 846.690 52.090 ;
        RECT 824.810 51.955 825.190 51.990 ;
        RECT 863.410 51.850 866.245 52.155 ;
        RECT 882.225 51.950 885.360 52.260 ;
        RECT 884.980 51.915 885.360 51.950 ;
        RECT 863.480 51.815 863.860 51.850 ;
        RECT 806.855 50.580 810.260 51.020 ;
        RECT 810.600 50.380 810.980 50.760 ;
        RECT 813.315 50.420 813.695 50.800 ;
        RECT 817.500 50.370 817.880 50.750 ;
        RECT 823.335 50.355 824.630 50.735 ;
        RECT 825.370 50.355 828.630 50.735 ;
        RECT 829.370 50.355 832.630 50.735 ;
        RECT 833.370 50.355 834.555 50.735 ;
        RECT 836.820 50.355 838.130 50.735 ;
        RECT 838.870 50.355 842.130 50.735 ;
        RECT 842.870 50.355 846.130 50.735 ;
        RECT 846.870 50.355 847.885 50.735 ;
        RECT 807.925 49.955 809.665 50.245 ;
        RECT 811.715 49.905 812.915 50.195 ;
        RECT 814.425 49.875 817.020 50.250 ;
        RECT 818.635 49.970 819.015 50.350 ;
        RECT 862.005 50.215 863.300 50.595 ;
        RECT 868.040 50.215 871.300 50.595 ;
        RECT 872.040 50.215 873.225 50.595 ;
        RECT 875.490 50.215 876.800 50.595 ;
        RECT 877.540 50.215 880.800 50.595 ;
        RECT 885.540 50.215 886.555 50.595 ;
        RECT 889.620 50.460 893.035 50.880 ;
        RECT 893.365 50.240 893.745 50.620 ;
        RECT 896.080 50.280 896.460 50.660 ;
        RECT 900.265 50.230 900.645 50.610 ;
        RECT 824.810 49.655 825.190 50.035 ;
        RECT 828.810 49.655 829.190 50.035 ;
        RECT 832.810 49.990 833.190 50.035 ;
        RECT 838.310 49.990 838.690 50.035 ;
        RECT 832.760 49.675 838.695 49.990 ;
        RECT 832.810 49.655 833.190 49.675 ;
        RECT 838.310 49.655 838.690 49.675 ;
        RECT 842.310 49.655 842.690 50.035 ;
        RECT 846.310 49.655 846.690 50.035 ;
        RECT 863.480 49.515 863.860 49.895 ;
        RECT 867.480 49.515 867.860 49.895 ;
        RECT 871.480 49.850 871.860 49.895 ;
        RECT 876.980 49.850 877.360 49.895 ;
        RECT 871.430 49.535 877.365 49.850 ;
        RECT 871.480 49.515 871.860 49.535 ;
        RECT 876.980 49.515 877.360 49.535 ;
        RECT 880.980 49.515 881.360 49.895 ;
        RECT 884.980 49.515 885.360 49.895 ;
        RECT 890.690 49.815 892.430 50.105 ;
        RECT 894.480 49.765 895.680 50.055 ;
        RECT 897.190 49.725 899.820 50.180 ;
        RECT 901.400 49.830 901.780 50.210 ;
        RECT 806.165 49.195 819.990 49.495 ;
        RECT 821.665 49.030 837.675 49.405 ;
        RECT 855.570 48.890 876.345 49.265 ;
        RECT 806.170 48.450 824.590 48.750 ;
        RECT 826.035 48.440 853.345 48.780 ;
        RECT 805.650 47.735 812.910 48.035 ;
        RECT 625.325 47.170 682.665 47.180 ;
        RECT 625.325 47.000 691.670 47.170 ;
        RECT 790.705 47.115 794.830 47.385 ;
        RECT 806.205 47.200 810.290 47.470 ;
        RECT 816.610 47.435 820.360 47.710 ;
        RECT 821.665 47.675 847.895 48.065 ;
        RECT 854.600 47.535 886.565 47.925 ;
        RECT 821.665 47.310 840.335 47.320 ;
        RECT 821.665 47.180 851.685 47.310 ;
        RECT 899.375 47.295 902.505 47.570 ;
        RECT 903.250 47.535 903.630 54.695 ;
        RECT 952.905 52.655 954.105 53.035 ;
        RECT 904.490 52.235 911.230 52.535 ;
        RECT 955.860 52.440 958.135 52.950 ;
        RECT 960.760 52.440 963.060 52.950 ;
        RECT 965.355 52.440 967.635 52.950 ;
        RECT 972.430 52.755 973.665 53.135 ;
        RECT 905.080 50.440 908.535 50.880 ;
        RECT 908.825 50.240 909.205 50.620 ;
        RECT 911.540 50.280 911.920 50.660 ;
        RECT 915.725 50.230 916.105 50.610 ;
        RECT 952.905 50.355 956.165 50.735 ;
        RECT 956.905 50.355 960.165 50.735 ;
        RECT 966.405 50.355 969.665 50.735 ;
        RECT 970.405 50.355 973.665 50.735 ;
        RECT 906.150 49.815 907.890 50.105 ;
        RECT 909.940 49.765 911.140 50.055 ;
        RECT 912.650 49.735 915.275 50.145 ;
        RECT 916.860 49.830 917.240 50.210 ;
        RECT 903.895 49.055 919.815 49.355 ;
        RECT 904.430 48.310 921.375 48.610 ;
        RECT 953.570 48.440 979.865 48.780 ;
        RECT 985.905 47.675 986.285 54.835 ;
        RECT 987.735 50.620 991.110 51.020 ;
        RECT 991.480 50.380 991.860 50.760 ;
        RECT 994.195 50.420 994.575 50.800 ;
        RECT 998.380 50.370 998.760 50.750 ;
        RECT 988.805 49.955 990.545 50.245 ;
        RECT 992.595 49.905 993.795 50.195 ;
        RECT 995.305 49.875 997.915 50.300 ;
        RECT 999.515 49.970 999.895 50.350 ;
        RECT 987.050 49.195 1000.615 49.510 ;
        RECT 987.045 48.450 1000.605 48.750 ;
        RECT 987.065 47.735 993.790 48.035 ;
        RECT 914.835 47.295 922.535 47.570 ;
        RECT 997.490 47.435 1000.595 47.710 ;
        RECT 1001.365 47.675 1001.745 54.835 ;
        RECT 1057.895 54.695 1114.250 54.835 ;
        RECT 1018.005 53.710 1055.555 53.850 ;
        RECT 1018.005 53.565 1083.655 53.710 ;
        RECT 1054.880 53.425 1083.655 53.565 ;
        RECT 1085.325 53.405 1092.030 53.705 ;
        RECT 1019.515 52.655 1020.970 53.035 ;
        RECT 1021.710 52.655 1022.910 53.035 ;
        RECT 1024.665 52.440 1026.940 52.950 ;
        RECT 1029.565 52.440 1031.865 52.950 ;
        RECT 1034.160 52.440 1036.440 52.950 ;
        RECT 1041.235 52.755 1042.470 53.135 ;
        RECT 1043.210 52.755 1044.490 53.135 ;
        RECT 1058.185 52.515 1059.640 52.895 ;
        RECT 1042.650 52.400 1043.030 52.435 ;
        RECT 1021.150 52.295 1021.530 52.335 ;
        RECT 1021.080 51.990 1023.915 52.295 ;
        RECT 1039.895 52.090 1043.030 52.400 ;
        RECT 1063.335 52.300 1065.610 52.810 ;
        RECT 1068.235 52.300 1070.535 52.810 ;
        RECT 1072.830 52.300 1075.110 52.810 ;
        RECT 1081.880 52.615 1083.160 52.995 ;
        RECT 1081.320 52.260 1081.700 52.295 ;
        RECT 1059.820 52.155 1060.200 52.195 ;
        RECT 1042.650 52.055 1043.030 52.090 ;
        RECT 1021.150 51.955 1021.530 51.990 ;
        RECT 1059.750 51.850 1062.585 52.155 ;
        RECT 1078.565 51.950 1081.700 52.260 ;
        RECT 1081.320 51.915 1081.700 51.950 ;
        RECT 1059.820 51.815 1060.200 51.850 ;
        RECT 1003.195 50.580 1006.600 51.020 ;
        RECT 1006.940 50.380 1007.320 50.760 ;
        RECT 1009.655 50.420 1010.035 50.800 ;
        RECT 1013.840 50.370 1014.220 50.750 ;
        RECT 1019.675 50.355 1020.970 50.735 ;
        RECT 1021.710 50.355 1024.970 50.735 ;
        RECT 1025.710 50.355 1028.970 50.735 ;
        RECT 1029.710 50.355 1030.895 50.735 ;
        RECT 1033.160 50.355 1034.470 50.735 ;
        RECT 1035.210 50.355 1038.470 50.735 ;
        RECT 1039.210 50.355 1042.470 50.735 ;
        RECT 1043.210 50.355 1044.225 50.735 ;
        RECT 1004.265 49.955 1006.005 50.245 ;
        RECT 1008.055 49.905 1009.255 50.195 ;
        RECT 1010.765 49.875 1013.360 50.250 ;
        RECT 1014.975 49.970 1015.355 50.350 ;
        RECT 1058.345 50.215 1059.640 50.595 ;
        RECT 1064.380 50.215 1067.640 50.595 ;
        RECT 1068.380 50.215 1069.565 50.595 ;
        RECT 1071.830 50.215 1073.140 50.595 ;
        RECT 1073.880 50.215 1077.140 50.595 ;
        RECT 1081.880 50.215 1082.895 50.595 ;
        RECT 1085.960 50.460 1089.375 50.880 ;
        RECT 1089.705 50.240 1090.085 50.620 ;
        RECT 1092.420 50.280 1092.800 50.660 ;
        RECT 1096.605 50.230 1096.985 50.610 ;
        RECT 1021.150 49.655 1021.530 50.035 ;
        RECT 1025.150 49.655 1025.530 50.035 ;
        RECT 1029.150 49.990 1029.530 50.035 ;
        RECT 1034.650 49.990 1035.030 50.035 ;
        RECT 1029.100 49.675 1035.035 49.990 ;
        RECT 1029.150 49.655 1029.530 49.675 ;
        RECT 1034.650 49.655 1035.030 49.675 ;
        RECT 1038.650 49.655 1039.030 50.035 ;
        RECT 1042.650 49.655 1043.030 50.035 ;
        RECT 1059.820 49.515 1060.200 49.895 ;
        RECT 1063.820 49.515 1064.200 49.895 ;
        RECT 1067.820 49.850 1068.200 49.895 ;
        RECT 1073.320 49.850 1073.700 49.895 ;
        RECT 1067.770 49.535 1073.705 49.850 ;
        RECT 1067.820 49.515 1068.200 49.535 ;
        RECT 1073.320 49.515 1073.700 49.535 ;
        RECT 1077.320 49.515 1077.700 49.895 ;
        RECT 1081.320 49.515 1081.700 49.895 ;
        RECT 1087.030 49.815 1088.770 50.105 ;
        RECT 1090.820 49.765 1092.020 50.055 ;
        RECT 1093.530 49.725 1096.160 50.180 ;
        RECT 1097.740 49.830 1098.120 50.210 ;
        RECT 1002.505 49.195 1016.330 49.495 ;
        RECT 1018.005 49.030 1034.015 49.405 ;
        RECT 1051.910 48.890 1072.685 49.265 ;
        RECT 1002.510 48.450 1020.930 48.750 ;
        RECT 1022.375 48.440 1049.685 48.780 ;
        RECT 1001.990 47.735 1009.250 48.035 ;
        RECT 821.665 47.170 879.005 47.180 ;
        RECT 821.665 47.000 888.010 47.170 ;
        RECT 987.045 47.115 991.170 47.385 ;
        RECT 1002.545 47.200 1006.630 47.470 ;
        RECT 1012.950 47.435 1016.700 47.710 ;
        RECT 1018.005 47.675 1044.235 48.065 ;
        RECT 1050.940 47.535 1082.905 47.925 ;
        RECT 1018.005 47.310 1036.675 47.320 ;
        RECT 1018.005 47.180 1048.025 47.310 ;
        RECT 1095.715 47.295 1098.845 47.570 ;
        RECT 1099.590 47.535 1099.970 54.695 ;
        RECT 1149.230 52.660 1150.430 53.040 ;
        RECT 1100.830 52.235 1107.570 52.535 ;
        RECT 1152.185 52.445 1154.460 52.955 ;
        RECT 1157.085 52.445 1159.385 52.955 ;
        RECT 1161.680 52.445 1163.960 52.955 ;
        RECT 1168.755 52.760 1169.990 53.140 ;
        RECT 1101.420 50.440 1104.875 50.880 ;
        RECT 1105.165 50.240 1105.545 50.620 ;
        RECT 1107.880 50.280 1108.260 50.660 ;
        RECT 1112.065 50.230 1112.445 50.610 ;
        RECT 1149.230 50.360 1152.490 50.740 ;
        RECT 1153.230 50.360 1156.490 50.740 ;
        RECT 1162.730 50.360 1165.990 50.740 ;
        RECT 1166.730 50.360 1169.990 50.740 ;
        RECT 1102.490 49.815 1104.230 50.105 ;
        RECT 1106.280 49.765 1107.480 50.055 ;
        RECT 1108.990 49.735 1111.615 50.145 ;
        RECT 1113.200 49.830 1113.580 50.210 ;
        RECT 1100.235 49.055 1116.155 49.355 ;
        RECT 1100.770 48.310 1117.715 48.610 ;
        RECT 1149.895 48.445 1176.190 48.785 ;
        RECT 1182.245 47.675 1182.625 54.835 ;
        RECT 1184.075 50.620 1187.450 51.020 ;
        RECT 1187.820 50.380 1188.200 50.760 ;
        RECT 1190.535 50.420 1190.915 50.800 ;
        RECT 1194.720 50.370 1195.100 50.750 ;
        RECT 1185.145 49.955 1186.885 50.245 ;
        RECT 1188.935 49.905 1190.135 50.195 ;
        RECT 1191.645 49.875 1194.255 50.300 ;
        RECT 1195.855 49.970 1196.235 50.350 ;
        RECT 1183.390 49.195 1196.955 49.510 ;
        RECT 1183.385 48.450 1196.945 48.750 ;
        RECT 1183.405 47.735 1190.130 48.035 ;
        RECT 1111.175 47.295 1118.875 47.570 ;
        RECT 1193.830 47.435 1196.935 47.710 ;
        RECT 1197.705 47.675 1198.085 54.835 ;
        RECT 1254.235 54.695 1310.590 54.835 ;
        RECT 1214.345 53.710 1251.895 53.850 ;
        RECT 1214.345 53.565 1279.995 53.710 ;
        RECT 1251.220 53.425 1279.995 53.565 ;
        RECT 1281.665 53.405 1288.370 53.705 ;
        RECT 1215.855 52.655 1217.310 53.035 ;
        RECT 1218.050 52.655 1219.250 53.035 ;
        RECT 1221.005 52.440 1223.280 52.950 ;
        RECT 1225.905 52.440 1228.205 52.950 ;
        RECT 1230.500 52.440 1232.780 52.950 ;
        RECT 1237.575 52.755 1238.810 53.135 ;
        RECT 1239.550 52.755 1240.830 53.135 ;
        RECT 1254.525 52.515 1255.980 52.895 ;
        RECT 1256.720 52.515 1257.920 52.895 ;
        RECT 1238.990 52.400 1239.370 52.435 ;
        RECT 1217.490 52.295 1217.870 52.335 ;
        RECT 1217.420 51.990 1220.255 52.295 ;
        RECT 1236.235 52.090 1239.370 52.400 ;
        RECT 1259.675 52.300 1261.950 52.810 ;
        RECT 1264.575 52.300 1266.875 52.810 ;
        RECT 1269.170 52.300 1271.450 52.810 ;
        RECT 1276.245 52.615 1277.480 52.995 ;
        RECT 1278.220 52.615 1279.500 52.995 ;
        RECT 1277.660 52.260 1278.040 52.295 ;
        RECT 1256.160 52.155 1256.540 52.195 ;
        RECT 1238.990 52.055 1239.370 52.090 ;
        RECT 1217.490 51.955 1217.870 51.990 ;
        RECT 1256.090 51.850 1258.925 52.155 ;
        RECT 1274.905 51.950 1278.040 52.260 ;
        RECT 1277.660 51.915 1278.040 51.950 ;
        RECT 1256.160 51.815 1256.540 51.850 ;
        RECT 1199.535 50.580 1202.940 51.020 ;
        RECT 1203.280 50.380 1203.660 50.760 ;
        RECT 1205.995 50.420 1206.375 50.800 ;
        RECT 1210.180 50.370 1210.560 50.750 ;
        RECT 1216.015 50.355 1217.310 50.735 ;
        RECT 1218.050 50.355 1221.310 50.735 ;
        RECT 1222.050 50.355 1225.310 50.735 ;
        RECT 1226.050 50.355 1227.235 50.735 ;
        RECT 1229.500 50.355 1230.810 50.735 ;
        RECT 1231.550 50.355 1234.810 50.735 ;
        RECT 1235.550 50.355 1238.810 50.735 ;
        RECT 1239.550 50.355 1240.565 50.735 ;
        RECT 1200.605 49.955 1202.345 50.245 ;
        RECT 1204.395 49.905 1205.595 50.195 ;
        RECT 1207.105 49.875 1209.700 50.250 ;
        RECT 1211.315 49.970 1211.695 50.350 ;
        RECT 1254.685 50.215 1255.980 50.595 ;
        RECT 1256.720 50.215 1259.980 50.595 ;
        RECT 1260.720 50.215 1263.980 50.595 ;
        RECT 1264.720 50.215 1265.905 50.595 ;
        RECT 1268.170 50.215 1269.480 50.595 ;
        RECT 1270.220 50.215 1273.480 50.595 ;
        RECT 1274.220 50.215 1277.480 50.595 ;
        RECT 1278.220 50.215 1279.235 50.595 ;
        RECT 1282.300 50.460 1285.715 50.880 ;
        RECT 1286.045 50.240 1286.425 50.620 ;
        RECT 1288.760 50.280 1289.140 50.660 ;
        RECT 1292.945 50.230 1293.325 50.610 ;
        RECT 1217.490 49.655 1217.870 50.035 ;
        RECT 1221.490 49.655 1221.870 50.035 ;
        RECT 1225.490 49.990 1225.870 50.035 ;
        RECT 1230.990 49.990 1231.370 50.035 ;
        RECT 1225.440 49.675 1231.375 49.990 ;
        RECT 1225.490 49.655 1225.870 49.675 ;
        RECT 1230.990 49.655 1231.370 49.675 ;
        RECT 1234.990 49.655 1235.370 50.035 ;
        RECT 1238.990 49.655 1239.370 50.035 ;
        RECT 1256.160 49.515 1256.540 49.895 ;
        RECT 1260.160 49.515 1260.540 49.895 ;
        RECT 1264.160 49.850 1264.540 49.895 ;
        RECT 1269.660 49.850 1270.040 49.895 ;
        RECT 1264.110 49.535 1270.045 49.850 ;
        RECT 1264.160 49.515 1264.540 49.535 ;
        RECT 1269.660 49.515 1270.040 49.535 ;
        RECT 1273.660 49.515 1274.040 49.895 ;
        RECT 1277.660 49.515 1278.040 49.895 ;
        RECT 1283.370 49.815 1285.110 50.105 ;
        RECT 1287.160 49.765 1288.360 50.055 ;
        RECT 1289.870 49.725 1292.500 50.180 ;
        RECT 1294.080 49.830 1294.460 50.210 ;
        RECT 1198.845 49.195 1212.670 49.495 ;
        RECT 1214.345 49.030 1230.355 49.405 ;
        RECT 1248.250 48.890 1269.025 49.265 ;
        RECT 1281.650 49.055 1295.265 49.355 ;
        RECT 1198.850 48.450 1217.270 48.750 ;
        RECT 1218.715 48.440 1246.025 48.780 ;
        RECT 1257.385 48.300 1279.940 48.640 ;
        RECT 1281.050 48.310 1295.695 48.610 ;
        RECT 1198.330 47.735 1205.590 48.035 ;
        RECT 1018.005 47.170 1075.345 47.180 ;
        RECT 1018.005 47.000 1084.350 47.170 ;
        RECT 1183.385 47.115 1187.510 47.385 ;
        RECT 1198.885 47.200 1202.970 47.470 ;
        RECT 1209.290 47.435 1213.040 47.710 ;
        RECT 1214.345 47.675 1240.575 48.065 ;
        RECT 1247.280 47.535 1279.245 47.925 ;
        RECT 1214.345 47.310 1233.015 47.320 ;
        RECT 1214.345 47.180 1244.365 47.310 ;
        RECT 1292.055 47.295 1295.185 47.570 ;
        RECT 1295.930 47.535 1296.310 54.695 ;
        RECT 1297.170 52.235 1303.910 52.535 ;
        RECT 1297.760 50.440 1301.215 50.880 ;
        RECT 1304.220 50.280 1304.600 50.660 ;
        RECT 1302.620 49.765 1303.820 50.055 ;
        RECT 1309.540 49.830 1309.920 50.210 ;
        RECT 1296.575 49.055 1312.495 49.355 ;
        RECT 1297.110 48.310 1314.055 48.610 ;
        RECT 1214.345 47.170 1271.685 47.180 ;
        RECT 1214.345 47.000 1280.690 47.170 ;
        RECT 6.460 46.555 10.590 46.855 ;
        RECT -59.665 45.735 -56.100 45.745 ;
        RECT -59.665 45.410 -55.305 45.735 ;
        RECT -9.340 45.490 -3.425 45.825 ;
        RECT -6.070 45.470 -3.425 45.490 ;
        RECT -56.260 45.400 -55.305 45.410 ;
        RECT -79.070 44.770 -75.770 45.150 ;
        RECT -75.070 44.770 -71.770 45.150 ;
        RECT -65.570 44.770 -62.270 45.150 ;
        RECT -61.570 44.770 -58.270 45.150 ;
        RECT -28.745 44.850 -25.445 45.230 ;
        RECT -24.745 44.850 -21.445 45.230 ;
        RECT -15.245 44.850 -11.945 45.230 ;
        RECT -11.245 44.850 -7.945 45.230 ;
        RECT -79.070 42.770 -77.785 43.150 ;
        RECT -59.755 42.770 -58.270 43.150 ;
        RECT -28.745 42.850 -27.460 43.230 ;
        RECT -9.430 42.850 -7.945 43.230 ;
        RECT -77.565 42.090 -76.045 42.450 ;
        RECT -27.240 42.170 -25.720 42.530 ;
        RECT 4.085 40.725 4.465 46.555 ;
        RECT 12.965 46.505 17.465 46.815 ;
        RECT 21.920 46.555 26.050 46.855 ;
        RECT 8.925 45.955 15.315 46.245 ;
        RECT 8.340 45.375 18.995 45.710 ;
        RECT 7.690 44.790 10.610 45.090 ;
        RECT 14.155 44.775 17.525 45.075 ;
        RECT 5.905 44.040 6.285 44.420 ;
        RECT 8.310 44.055 10.090 44.345 ;
        RECT 11.565 44.145 12.755 44.430 ;
        RECT 15.685 44.025 16.995 44.345 ;
        RECT 7.040 43.440 7.420 43.820 ;
        RECT 10.785 43.480 11.165 43.860 ;
        RECT 13.495 43.470 13.875 43.850 ;
        RECT 14.905 43.315 18.085 43.635 ;
        RECT 4.835 40.725 8.930 40.730 ;
        RECT 19.545 40.725 19.925 46.555 ;
        RECT 28.425 46.505 32.925 46.815 ;
        RECT 120.145 46.415 124.275 46.715 ;
        RECT 24.385 45.955 30.775 46.245 ;
        RECT 35.655 46.205 71.565 46.345 ;
        RECT 35.655 46.075 102.930 46.205 ;
        RECT 71.185 45.935 102.930 46.075 ;
        RECT 23.800 45.375 34.305 45.710 ;
        RECT 59.275 45.510 69.825 45.845 ;
        RECT 107.150 45.815 113.540 46.105 ;
        RECT 23.150 44.790 26.070 45.090 ;
        RECT 29.615 44.775 32.985 45.075 ;
        RECT 37.865 44.870 39.170 45.250 ;
        RECT 39.870 44.870 43.170 45.250 ;
        RECT 43.870 44.870 47.170 45.250 ;
        RECT 47.870 44.870 49.230 45.250 ;
        RECT 51.205 44.870 52.670 45.250 ;
        RECT 53.370 44.870 56.670 45.250 ;
        RECT 57.370 44.870 60.670 45.250 ;
        RECT 61.370 44.870 62.550 45.250 ;
        RECT 106.565 45.235 117.045 45.570 ;
        RECT 76.535 44.730 77.840 45.110 ;
        RECT 82.540 44.730 85.840 45.110 ;
        RECT 86.540 44.730 87.900 45.110 ;
        RECT 89.875 44.730 91.340 45.110 ;
        RECT 92.040 44.730 95.340 45.110 ;
        RECT 100.040 44.730 101.220 45.110 ;
        RECT 39.330 44.525 39.710 44.560 ;
        RECT 21.365 44.040 21.745 44.420 ;
        RECT 23.770 44.055 25.550 44.345 ;
        RECT 27.025 44.145 28.215 44.430 ;
        RECT 31.145 44.025 32.455 44.345 ;
        RECT 39.065 44.215 42.075 44.525 ;
        RECT 39.330 44.180 39.710 44.215 ;
        RECT 43.330 44.180 44.420 44.560 ;
        RECT 47.330 44.555 47.710 44.560 ;
        RECT 44.850 44.190 47.715 44.555 ;
        RECT 52.830 44.535 53.210 44.560 ;
        RECT 52.815 44.215 54.960 44.535 ;
        RECT 47.330 44.180 47.710 44.190 ;
        RECT 52.830 44.180 53.210 44.215 ;
        RECT 55.875 44.180 57.210 44.560 ;
        RECT 60.830 44.540 61.210 44.560 ;
        RECT 58.365 44.220 61.275 44.540 ;
        RECT 78.000 44.385 78.380 44.420 ;
        RECT 60.830 44.180 61.210 44.220 ;
        RECT 77.735 44.075 80.745 44.385 ;
        RECT 78.000 44.040 78.380 44.075 ;
        RECT 82.000 44.040 83.090 44.420 ;
        RECT 86.000 44.415 86.380 44.420 ;
        RECT 83.520 44.050 86.385 44.415 ;
        RECT 91.500 44.395 91.880 44.420 ;
        RECT 91.485 44.075 93.630 44.395 ;
        RECT 86.000 44.040 86.380 44.050 ;
        RECT 91.500 44.040 91.880 44.075 ;
        RECT 94.545 44.040 95.880 44.420 ;
        RECT 99.500 44.400 99.880 44.420 ;
        RECT 97.035 44.080 99.945 44.400 ;
        RECT 99.500 44.040 99.880 44.080 ;
        RECT 104.130 43.900 104.510 44.280 ;
        RECT 106.535 43.915 108.315 44.205 ;
        RECT 109.790 44.005 110.980 44.290 ;
        RECT 113.910 43.885 115.220 44.205 ;
        RECT 22.500 43.440 22.880 43.820 ;
        RECT 26.245 43.480 26.625 43.860 ;
        RECT 28.955 43.470 29.335 43.850 ;
        RECT 30.365 43.315 33.545 43.635 ;
        RECT 105.265 43.300 105.645 43.680 ;
        RECT 109.010 43.340 109.390 43.720 ;
        RECT 111.720 43.330 112.100 43.710 ;
        RECT 37.680 42.870 39.170 43.250 ;
        RECT 39.870 42.870 41.155 43.250 ;
        RECT 59.185 42.870 60.670 43.250 ;
        RECT 61.370 42.870 62.445 43.250 ;
        RECT 113.130 43.175 116.310 43.495 ;
        RECT 76.350 42.730 77.840 43.110 ;
        RECT 100.040 42.730 101.115 43.110 ;
        RECT 39.330 42.180 40.420 42.560 ;
        RECT 41.375 42.190 42.895 42.550 ;
        RECT 43.815 42.185 56.665 42.520 ;
        RECT 60.830 42.515 61.210 42.560 ;
        RECT 60.095 42.215 61.405 42.515 ;
        RECT 60.830 42.180 61.210 42.215 ;
        RECT 78.000 42.040 79.090 42.420 ;
        RECT 80.045 42.050 81.565 42.410 ;
        RECT 82.485 42.045 95.335 42.380 ;
        RECT 99.500 42.375 99.880 42.420 ;
        RECT 98.765 42.075 100.075 42.375 ;
        RECT 99.500 42.040 99.880 42.075 ;
        RECT 36.185 41.545 69.265 41.670 ;
        RECT 36.185 41.320 101.510 41.545 ;
        RECT 68.560 41.180 101.510 41.320 ;
        RECT 103.305 41.170 107.565 41.525 ;
        RECT 20.295 40.725 24.390 40.730 ;
        RECT 3.715 40.720 8.930 40.725 ;
        RECT 19.175 40.720 24.390 40.725 ;
        RECT 34.635 40.720 74.885 40.725 ;
        RECT -82.755 39.725 -56.100 40.625 ;
        RECT -32.430 39.805 -5.775 40.705 ;
        RECT 3.715 40.585 74.885 40.720 ;
        RECT 101.510 40.585 107.155 40.590 ;
        RECT 117.770 40.585 118.150 46.415 ;
        RECT 126.650 46.365 131.150 46.675 ;
        RECT 202.825 46.555 206.955 46.855 ;
        RECT 122.610 45.815 129.000 46.105 ;
        RECT 122.025 45.235 138.045 45.570 ;
        RECT 186.830 45.500 192.745 45.835 ;
        RECT 190.100 45.480 192.745 45.500 ;
        RECT 121.375 44.650 124.295 44.950 ;
        RECT 127.840 44.635 131.210 44.935 ;
        RECT 167.425 44.860 170.725 45.240 ;
        RECT 171.425 44.860 174.725 45.240 ;
        RECT 180.925 44.860 184.225 45.240 ;
        RECT 184.925 44.860 188.225 45.240 ;
        RECT 119.590 43.900 119.970 44.280 ;
        RECT 121.995 43.915 123.775 44.205 ;
        RECT 125.250 44.005 126.440 44.290 ;
        RECT 129.370 43.885 130.680 44.205 ;
        RECT 120.725 43.300 121.105 43.680 ;
        RECT 124.470 43.340 124.850 43.720 ;
        RECT 127.180 43.330 127.560 43.710 ;
        RECT 128.590 43.175 131.770 43.495 ;
        RECT 167.425 42.860 168.710 43.240 ;
        RECT 186.740 42.860 188.225 43.240 ;
        RECT 118.870 42.090 123.020 42.360 ;
        RECT 168.930 42.180 170.450 42.540 ;
        RECT 200.450 40.725 200.830 46.555 ;
        RECT 209.330 46.505 213.830 46.815 ;
        RECT 218.285 46.555 222.415 46.855 ;
        RECT 458.730 46.825 495.295 46.965 ;
        RECT 655.105 46.860 691.670 47.000 ;
        RECT 851.445 46.860 888.010 47.000 ;
        RECT 1047.785 46.860 1084.350 47.000 ;
        RECT 1244.125 46.860 1280.690 47.000 ;
        RECT 205.290 45.955 211.680 46.245 ;
        RECT 204.705 45.375 215.360 45.710 ;
        RECT 204.055 44.790 206.975 45.090 ;
        RECT 210.520 44.775 213.890 45.075 ;
        RECT 202.270 44.040 202.650 44.420 ;
        RECT 204.675 44.055 206.455 44.345 ;
        RECT 207.930 44.145 209.120 44.430 ;
        RECT 212.050 44.025 213.360 44.345 ;
        RECT 203.405 43.440 203.785 43.820 ;
        RECT 207.150 43.480 207.530 43.860 ;
        RECT 209.860 43.470 210.240 43.850 ;
        RECT 211.270 43.315 214.450 43.635 ;
        RECT 201.200 40.725 205.295 40.730 ;
        RECT 215.910 40.725 216.290 46.555 ;
        RECT 224.790 46.505 229.290 46.815 ;
        RECT 316.510 46.415 320.640 46.715 ;
        RECT 220.750 45.955 227.140 46.245 ;
        RECT 232.020 46.205 267.930 46.345 ;
        RECT 232.020 46.075 299.295 46.205 ;
        RECT 267.550 45.935 299.295 46.075 ;
        RECT 220.165 45.375 230.670 45.710 ;
        RECT 255.640 45.510 266.190 45.845 ;
        RECT 303.515 45.815 309.905 46.105 ;
        RECT 219.515 44.790 222.435 45.090 ;
        RECT 225.980 44.775 229.350 45.075 ;
        RECT 234.230 44.870 235.535 45.250 ;
        RECT 236.235 44.870 239.535 45.250 ;
        RECT 240.235 44.870 243.535 45.250 ;
        RECT 244.235 44.870 245.595 45.250 ;
        RECT 247.570 44.870 249.035 45.250 ;
        RECT 249.735 44.870 253.035 45.250 ;
        RECT 253.735 44.870 257.035 45.250 ;
        RECT 257.735 44.870 258.915 45.250 ;
        RECT 302.930 45.235 313.410 45.570 ;
        RECT 272.900 44.730 274.205 45.110 ;
        RECT 278.905 44.730 282.205 45.110 ;
        RECT 282.905 44.730 284.265 45.110 ;
        RECT 286.240 44.730 287.705 45.110 ;
        RECT 288.405 44.730 291.705 45.110 ;
        RECT 296.405 44.730 297.585 45.110 ;
        RECT 235.695 44.525 236.075 44.560 ;
        RECT 217.730 44.040 218.110 44.420 ;
        RECT 220.135 44.055 221.915 44.345 ;
        RECT 223.390 44.145 224.580 44.430 ;
        RECT 227.510 44.025 228.820 44.345 ;
        RECT 235.430 44.215 238.440 44.525 ;
        RECT 235.695 44.180 236.075 44.215 ;
        RECT 239.695 44.180 240.785 44.560 ;
        RECT 243.695 44.555 244.075 44.560 ;
        RECT 241.215 44.190 244.080 44.555 ;
        RECT 249.195 44.535 249.575 44.560 ;
        RECT 249.180 44.215 251.325 44.535 ;
        RECT 243.695 44.180 244.075 44.190 ;
        RECT 249.195 44.180 249.575 44.215 ;
        RECT 252.240 44.180 253.575 44.560 ;
        RECT 257.195 44.540 257.575 44.560 ;
        RECT 254.730 44.220 257.640 44.540 ;
        RECT 274.365 44.385 274.745 44.420 ;
        RECT 257.195 44.180 257.575 44.220 ;
        RECT 274.100 44.075 277.110 44.385 ;
        RECT 274.365 44.040 274.745 44.075 ;
        RECT 278.365 44.040 279.455 44.420 ;
        RECT 282.365 44.415 282.745 44.420 ;
        RECT 279.885 44.050 282.750 44.415 ;
        RECT 287.865 44.395 288.245 44.420 ;
        RECT 287.850 44.075 289.995 44.395 ;
        RECT 282.365 44.040 282.745 44.050 ;
        RECT 287.865 44.040 288.245 44.075 ;
        RECT 290.910 44.040 292.245 44.420 ;
        RECT 295.865 44.400 296.245 44.420 ;
        RECT 293.400 44.080 296.310 44.400 ;
        RECT 295.865 44.040 296.245 44.080 ;
        RECT 300.495 43.900 300.875 44.280 ;
        RECT 302.900 43.915 304.680 44.205 ;
        RECT 306.155 44.005 307.345 44.290 ;
        RECT 310.275 43.885 311.585 44.205 ;
        RECT 218.865 43.440 219.245 43.820 ;
        RECT 222.610 43.480 222.990 43.860 ;
        RECT 225.320 43.470 225.700 43.850 ;
        RECT 226.730 43.315 229.910 43.635 ;
        RECT 301.630 43.300 302.010 43.680 ;
        RECT 305.375 43.340 305.755 43.720 ;
        RECT 308.085 43.330 308.465 43.710 ;
        RECT 234.045 42.870 235.535 43.250 ;
        RECT 236.235 42.870 237.520 43.250 ;
        RECT 255.550 42.870 257.035 43.250 ;
        RECT 257.735 42.870 258.810 43.250 ;
        RECT 309.495 43.175 312.675 43.495 ;
        RECT 272.715 42.730 274.205 43.110 ;
        RECT 296.405 42.730 297.480 43.110 ;
        RECT 235.695 42.180 236.785 42.560 ;
        RECT 237.740 42.190 239.260 42.550 ;
        RECT 240.180 42.185 253.030 42.520 ;
        RECT 257.195 42.515 257.575 42.560 ;
        RECT 256.460 42.215 257.770 42.515 ;
        RECT 257.195 42.180 257.575 42.215 ;
        RECT 274.365 42.040 275.455 42.420 ;
        RECT 276.410 42.050 277.930 42.410 ;
        RECT 278.850 42.045 291.700 42.380 ;
        RECT 295.865 42.375 296.245 42.420 ;
        RECT 295.130 42.075 296.440 42.375 ;
        RECT 295.865 42.040 296.245 42.075 ;
        RECT 232.550 41.545 265.630 41.670 ;
        RECT 232.550 41.320 297.875 41.545 ;
        RECT 264.925 41.180 297.875 41.320 ;
        RECT 299.670 41.170 303.930 41.525 ;
        RECT 216.660 40.725 220.755 40.730 ;
        RECT 200.080 40.720 205.295 40.725 ;
        RECT 215.540 40.720 220.755 40.725 ;
        RECT 231.000 40.720 271.250 40.725 ;
        RECT 118.520 40.585 122.615 40.590 ;
        RECT 3.715 40.580 107.155 40.585 ;
        RECT 117.400 40.580 122.615 40.585 ;
        RECT 3.715 39.825 132.430 40.580 ;
        RECT 74.855 39.685 132.430 39.825 ;
        RECT 163.740 39.815 190.395 40.715 ;
        RECT 200.080 40.585 271.250 40.720 ;
        RECT 297.875 40.585 303.520 40.590 ;
        RECT 314.135 40.585 314.515 46.415 ;
        RECT 323.015 46.365 327.515 46.675 ;
        RECT 399.225 46.505 403.355 46.805 ;
        RECT 318.975 45.815 325.365 46.105 ;
        RECT 318.390 45.235 334.410 45.570 ;
        RECT 383.220 45.460 389.135 45.795 ;
        RECT 386.490 45.440 389.135 45.460 ;
        RECT 317.740 44.650 320.660 44.950 ;
        RECT 324.205 44.635 327.575 44.935 ;
        RECT 363.815 44.820 367.115 45.200 ;
        RECT 367.815 44.820 371.115 45.200 ;
        RECT 377.315 44.820 380.615 45.200 ;
        RECT 381.315 44.820 384.615 45.200 ;
        RECT 315.955 43.900 316.335 44.280 ;
        RECT 318.360 43.915 320.140 44.205 ;
        RECT 321.615 44.005 322.805 44.290 ;
        RECT 325.735 43.885 327.045 44.205 ;
        RECT 317.090 43.300 317.470 43.680 ;
        RECT 320.835 43.340 321.215 43.720 ;
        RECT 323.545 43.330 323.925 43.710 ;
        RECT 324.955 43.175 328.135 43.495 ;
        RECT 363.815 42.820 365.100 43.200 ;
        RECT 383.130 42.820 384.615 43.200 ;
        RECT 315.235 42.090 319.385 42.360 ;
        RECT 365.320 42.140 366.840 42.500 ;
        RECT 396.850 40.675 397.230 46.505 ;
        RECT 405.730 46.455 410.230 46.765 ;
        RECT 414.685 46.505 418.815 46.805 ;
        RECT 401.690 45.905 408.080 46.195 ;
        RECT 401.105 45.325 411.760 45.660 ;
        RECT 400.455 44.740 403.375 45.040 ;
        RECT 406.920 44.725 410.290 45.025 ;
        RECT 398.670 43.990 399.050 44.370 ;
        RECT 401.075 44.005 402.855 44.295 ;
        RECT 404.330 44.095 405.520 44.380 ;
        RECT 408.450 43.975 409.760 44.295 ;
        RECT 399.805 43.390 400.185 43.770 ;
        RECT 403.550 43.430 403.930 43.810 ;
        RECT 406.260 43.420 406.640 43.800 ;
        RECT 407.670 43.265 410.850 43.585 ;
        RECT 397.600 40.675 401.695 40.680 ;
        RECT 412.310 40.675 412.690 46.505 ;
        RECT 421.190 46.455 425.690 46.765 ;
        RECT 512.910 46.365 517.040 46.665 ;
        RECT 417.150 45.905 423.540 46.195 ;
        RECT 428.420 46.155 464.330 46.295 ;
        RECT 428.420 46.025 495.695 46.155 ;
        RECT 463.950 45.885 495.695 46.025 ;
        RECT 416.565 45.325 427.070 45.660 ;
        RECT 452.040 45.460 462.590 45.795 ;
        RECT 499.915 45.765 506.305 46.055 ;
        RECT 415.915 44.740 418.835 45.040 ;
        RECT 422.380 44.725 425.750 45.025 ;
        RECT 430.630 44.820 431.935 45.200 ;
        RECT 432.635 44.820 435.935 45.200 ;
        RECT 436.635 44.820 439.935 45.200 ;
        RECT 440.635 44.820 441.995 45.200 ;
        RECT 443.970 44.820 445.435 45.200 ;
        RECT 446.135 44.820 449.435 45.200 ;
        RECT 450.135 44.820 453.435 45.200 ;
        RECT 454.135 44.820 455.315 45.200 ;
        RECT 499.330 45.185 509.810 45.520 ;
        RECT 469.300 44.680 470.605 45.060 ;
        RECT 475.305 44.680 478.605 45.060 ;
        RECT 479.305 44.680 480.665 45.060 ;
        RECT 482.640 44.680 484.105 45.060 ;
        RECT 484.805 44.680 488.105 45.060 ;
        RECT 492.805 44.680 493.985 45.060 ;
        RECT 432.095 44.475 432.475 44.510 ;
        RECT 414.130 43.990 414.510 44.370 ;
        RECT 416.535 44.005 418.315 44.295 ;
        RECT 419.790 44.095 420.980 44.380 ;
        RECT 423.910 43.975 425.220 44.295 ;
        RECT 431.830 44.165 434.840 44.475 ;
        RECT 432.095 44.130 432.475 44.165 ;
        RECT 436.095 44.130 437.185 44.510 ;
        RECT 440.095 44.505 440.475 44.510 ;
        RECT 437.615 44.140 440.480 44.505 ;
        RECT 445.595 44.485 445.975 44.510 ;
        RECT 445.580 44.165 447.725 44.485 ;
        RECT 440.095 44.130 440.475 44.140 ;
        RECT 445.595 44.130 445.975 44.165 ;
        RECT 448.640 44.130 449.975 44.510 ;
        RECT 453.595 44.490 453.975 44.510 ;
        RECT 451.130 44.170 454.040 44.490 ;
        RECT 470.765 44.335 471.145 44.370 ;
        RECT 453.595 44.130 453.975 44.170 ;
        RECT 470.500 44.025 473.510 44.335 ;
        RECT 470.765 43.990 471.145 44.025 ;
        RECT 474.765 43.990 475.855 44.370 ;
        RECT 478.765 44.365 479.145 44.370 ;
        RECT 476.285 44.000 479.150 44.365 ;
        RECT 484.265 44.345 484.645 44.370 ;
        RECT 484.250 44.025 486.395 44.345 ;
        RECT 478.765 43.990 479.145 44.000 ;
        RECT 484.265 43.990 484.645 44.025 ;
        RECT 487.310 43.990 488.645 44.370 ;
        RECT 492.265 44.350 492.645 44.370 ;
        RECT 489.800 44.030 492.710 44.350 ;
        RECT 492.265 43.990 492.645 44.030 ;
        RECT 496.895 43.850 497.275 44.230 ;
        RECT 499.300 43.865 501.080 44.155 ;
        RECT 502.555 43.955 503.745 44.240 ;
        RECT 506.675 43.835 507.985 44.155 ;
        RECT 415.265 43.390 415.645 43.770 ;
        RECT 419.010 43.430 419.390 43.810 ;
        RECT 421.720 43.420 422.100 43.800 ;
        RECT 423.130 43.265 426.310 43.585 ;
        RECT 498.030 43.250 498.410 43.630 ;
        RECT 501.775 43.290 502.155 43.670 ;
        RECT 504.485 43.280 504.865 43.660 ;
        RECT 430.445 42.820 431.935 43.200 ;
        RECT 432.635 42.820 433.920 43.200 ;
        RECT 451.950 42.820 453.435 43.200 ;
        RECT 454.135 42.820 455.210 43.200 ;
        RECT 505.895 43.125 509.075 43.445 ;
        RECT 469.115 42.680 470.605 43.060 ;
        RECT 492.805 42.680 493.880 43.060 ;
        RECT 432.095 42.130 433.185 42.510 ;
        RECT 434.140 42.140 435.660 42.500 ;
        RECT 436.580 42.135 449.430 42.470 ;
        RECT 453.595 42.465 453.975 42.510 ;
        RECT 452.860 42.165 454.170 42.465 ;
        RECT 453.595 42.130 453.975 42.165 ;
        RECT 470.765 41.990 471.855 42.370 ;
        RECT 472.810 42.000 474.330 42.360 ;
        RECT 475.250 41.995 488.100 42.330 ;
        RECT 492.265 42.325 492.645 42.370 ;
        RECT 491.530 42.025 492.840 42.325 ;
        RECT 492.265 41.990 492.645 42.025 ;
        RECT 428.950 41.495 462.030 41.620 ;
        RECT 428.950 41.270 494.275 41.495 ;
        RECT 461.325 41.130 494.275 41.270 ;
        RECT 496.070 41.120 500.330 41.475 ;
        RECT 413.060 40.675 417.155 40.680 ;
        RECT 314.885 40.585 318.980 40.590 ;
        RECT 200.080 40.580 303.520 40.585 ;
        RECT 313.765 40.580 318.980 40.585 ;
        RECT 200.080 39.825 328.795 40.580 ;
        RECT 271.220 39.685 328.795 39.825 ;
        RECT 360.130 39.775 386.785 40.675 ;
        RECT 396.480 40.670 401.695 40.675 ;
        RECT 411.940 40.670 417.155 40.675 ;
        RECT 427.400 40.670 467.650 40.675 ;
        RECT 396.480 40.535 467.650 40.670 ;
        RECT 494.275 40.535 499.920 40.540 ;
        RECT 510.535 40.535 510.915 46.365 ;
        RECT 519.415 46.315 523.915 46.625 ;
        RECT 595.600 46.540 599.730 46.840 ;
        RECT 515.375 45.765 521.765 46.055 ;
        RECT 514.790 45.185 530.810 45.520 ;
        RECT 579.540 45.505 585.455 45.840 ;
        RECT 582.810 45.485 585.455 45.505 ;
        RECT 514.140 44.600 517.060 44.900 ;
        RECT 520.605 44.585 523.975 44.885 ;
        RECT 560.135 44.865 563.435 45.245 ;
        RECT 564.135 44.865 567.435 45.245 ;
        RECT 573.635 44.865 576.935 45.245 ;
        RECT 577.635 44.865 580.935 45.245 ;
        RECT 512.355 43.850 512.735 44.230 ;
        RECT 514.760 43.865 516.540 44.155 ;
        RECT 518.015 43.955 519.205 44.240 ;
        RECT 522.135 43.835 523.445 44.155 ;
        RECT 513.490 43.250 513.870 43.630 ;
        RECT 517.235 43.290 517.615 43.670 ;
        RECT 519.945 43.280 520.325 43.660 ;
        RECT 521.355 43.125 524.535 43.445 ;
        RECT 560.135 42.865 561.420 43.245 ;
        RECT 579.450 42.865 580.935 43.245 ;
        RECT 511.635 42.040 515.785 42.310 ;
        RECT 561.640 42.185 563.160 42.545 ;
        RECT 511.285 40.535 515.380 40.540 ;
        RECT 396.480 40.530 499.920 40.535 ;
        RECT 510.165 40.530 515.380 40.535 ;
        RECT 396.480 39.775 525.195 40.530 ;
        RECT 556.450 39.820 583.105 40.720 ;
        RECT 593.225 40.710 593.605 46.540 ;
        RECT 602.105 46.490 606.605 46.800 ;
        RECT 611.060 46.540 615.190 46.840 ;
        RECT 598.065 45.940 604.455 46.230 ;
        RECT 597.480 45.360 608.135 45.695 ;
        RECT 596.830 44.775 599.750 45.075 ;
        RECT 603.295 44.760 606.665 45.060 ;
        RECT 595.045 44.025 595.425 44.405 ;
        RECT 597.450 44.040 599.230 44.330 ;
        RECT 600.705 44.130 601.895 44.415 ;
        RECT 604.825 44.010 606.135 44.330 ;
        RECT 596.180 43.425 596.560 43.805 ;
        RECT 599.925 43.465 600.305 43.845 ;
        RECT 602.635 43.455 603.015 43.835 ;
        RECT 604.045 43.300 607.225 43.620 ;
        RECT 593.975 40.710 598.070 40.715 ;
        RECT 608.685 40.710 609.065 46.540 ;
        RECT 617.565 46.490 622.065 46.800 ;
        RECT 709.285 46.400 713.415 46.700 ;
        RECT 613.525 45.940 619.915 46.230 ;
        RECT 624.795 46.190 660.705 46.330 ;
        RECT 624.795 46.060 692.070 46.190 ;
        RECT 660.325 45.920 692.070 46.060 ;
        RECT 612.940 45.360 623.445 45.695 ;
        RECT 648.415 45.495 658.965 45.830 ;
        RECT 696.290 45.800 702.680 46.090 ;
        RECT 612.290 44.775 615.210 45.075 ;
        RECT 618.755 44.760 622.125 45.060 ;
        RECT 627.005 44.855 628.310 45.235 ;
        RECT 629.010 44.855 632.310 45.235 ;
        RECT 633.010 44.855 636.310 45.235 ;
        RECT 637.010 44.855 638.370 45.235 ;
        RECT 640.345 44.855 641.810 45.235 ;
        RECT 642.510 44.855 645.810 45.235 ;
        RECT 646.510 44.855 649.810 45.235 ;
        RECT 650.510 44.855 651.690 45.235 ;
        RECT 695.705 45.220 706.185 45.555 ;
        RECT 665.675 44.715 666.980 45.095 ;
        RECT 671.680 44.715 674.980 45.095 ;
        RECT 675.680 44.715 677.040 45.095 ;
        RECT 679.015 44.715 680.480 45.095 ;
        RECT 681.180 44.715 684.480 45.095 ;
        RECT 689.180 44.715 690.360 45.095 ;
        RECT 628.470 44.510 628.850 44.545 ;
        RECT 610.505 44.025 610.885 44.405 ;
        RECT 612.910 44.040 614.690 44.330 ;
        RECT 616.165 44.130 617.355 44.415 ;
        RECT 620.285 44.010 621.595 44.330 ;
        RECT 628.205 44.200 631.215 44.510 ;
        RECT 628.470 44.165 628.850 44.200 ;
        RECT 632.470 44.165 633.560 44.545 ;
        RECT 636.470 44.540 636.850 44.545 ;
        RECT 633.990 44.175 636.855 44.540 ;
        RECT 641.970 44.520 642.350 44.545 ;
        RECT 641.955 44.200 644.100 44.520 ;
        RECT 636.470 44.165 636.850 44.175 ;
        RECT 641.970 44.165 642.350 44.200 ;
        RECT 645.015 44.165 646.350 44.545 ;
        RECT 649.970 44.525 650.350 44.545 ;
        RECT 647.505 44.205 650.415 44.525 ;
        RECT 667.140 44.370 667.520 44.405 ;
        RECT 649.970 44.165 650.350 44.205 ;
        RECT 666.875 44.060 669.885 44.370 ;
        RECT 667.140 44.025 667.520 44.060 ;
        RECT 671.140 44.025 672.230 44.405 ;
        RECT 675.140 44.400 675.520 44.405 ;
        RECT 672.660 44.035 675.525 44.400 ;
        RECT 680.640 44.380 681.020 44.405 ;
        RECT 680.625 44.060 682.770 44.380 ;
        RECT 675.140 44.025 675.520 44.035 ;
        RECT 680.640 44.025 681.020 44.060 ;
        RECT 683.685 44.025 685.020 44.405 ;
        RECT 688.640 44.385 689.020 44.405 ;
        RECT 686.175 44.065 689.085 44.385 ;
        RECT 688.640 44.025 689.020 44.065 ;
        RECT 693.270 43.885 693.650 44.265 ;
        RECT 695.675 43.900 697.455 44.190 ;
        RECT 698.930 43.990 700.120 44.275 ;
        RECT 703.050 43.870 704.360 44.190 ;
        RECT 611.640 43.425 612.020 43.805 ;
        RECT 615.385 43.465 615.765 43.845 ;
        RECT 618.095 43.455 618.475 43.835 ;
        RECT 619.505 43.300 622.685 43.620 ;
        RECT 694.405 43.285 694.785 43.665 ;
        RECT 698.150 43.325 698.530 43.705 ;
        RECT 700.860 43.315 701.240 43.695 ;
        RECT 626.820 42.855 628.310 43.235 ;
        RECT 629.010 42.855 630.295 43.235 ;
        RECT 648.325 42.855 649.810 43.235 ;
        RECT 650.510 42.855 651.585 43.235 ;
        RECT 702.270 43.160 705.450 43.480 ;
        RECT 665.490 42.715 666.980 43.095 ;
        RECT 689.180 42.715 690.255 43.095 ;
        RECT 628.470 42.165 629.560 42.545 ;
        RECT 630.515 42.175 632.035 42.535 ;
        RECT 632.955 42.170 645.805 42.505 ;
        RECT 649.970 42.500 650.350 42.545 ;
        RECT 649.235 42.200 650.545 42.500 ;
        RECT 649.970 42.165 650.350 42.200 ;
        RECT 667.140 42.025 668.230 42.405 ;
        RECT 669.185 42.035 670.705 42.395 ;
        RECT 671.625 42.030 684.475 42.365 ;
        RECT 688.640 42.360 689.020 42.405 ;
        RECT 687.905 42.060 689.215 42.360 ;
        RECT 688.640 42.025 689.020 42.060 ;
        RECT 625.325 41.530 658.405 41.655 ;
        RECT 625.325 41.305 690.650 41.530 ;
        RECT 657.700 41.165 690.650 41.305 ;
        RECT 692.445 41.155 696.705 41.510 ;
        RECT 609.435 40.710 613.530 40.715 ;
        RECT 592.855 40.705 598.070 40.710 ;
        RECT 608.315 40.705 613.530 40.710 ;
        RECT 623.775 40.705 664.025 40.710 ;
        RECT 592.855 40.570 664.025 40.705 ;
        RECT 690.650 40.570 696.295 40.575 ;
        RECT 706.910 40.570 707.290 46.400 ;
        RECT 715.790 46.350 720.290 46.660 ;
        RECT 791.940 46.540 796.070 46.840 ;
        RECT 711.750 45.800 718.140 46.090 ;
        RECT 711.165 45.220 727.185 45.555 ;
        RECT 775.905 45.510 781.820 45.845 ;
        RECT 779.175 45.490 781.820 45.510 ;
        RECT 710.515 44.635 713.435 44.935 ;
        RECT 716.980 44.620 720.350 44.920 ;
        RECT 756.500 44.870 759.800 45.250 ;
        RECT 760.500 44.870 763.800 45.250 ;
        RECT 770.000 44.870 773.300 45.250 ;
        RECT 774.000 44.870 777.300 45.250 ;
        RECT 708.730 43.885 709.110 44.265 ;
        RECT 711.135 43.900 712.915 44.190 ;
        RECT 714.390 43.990 715.580 44.275 ;
        RECT 718.510 43.870 719.820 44.190 ;
        RECT 709.865 43.285 710.245 43.665 ;
        RECT 713.610 43.325 713.990 43.705 ;
        RECT 716.320 43.315 716.700 43.695 ;
        RECT 717.730 43.160 720.910 43.480 ;
        RECT 756.500 42.870 757.785 43.250 ;
        RECT 775.815 42.870 777.300 43.250 ;
        RECT 708.010 42.075 712.160 42.345 ;
        RECT 758.005 42.190 759.525 42.550 ;
        RECT 707.660 40.570 711.755 40.575 ;
        RECT 592.855 40.565 696.295 40.570 ;
        RECT 706.540 40.565 711.755 40.570 ;
        RECT 592.855 39.810 721.570 40.565 ;
        RECT 752.815 39.825 779.470 40.725 ;
        RECT 789.565 40.710 789.945 46.540 ;
        RECT 798.445 46.490 802.945 46.800 ;
        RECT 807.400 46.540 811.530 46.840 ;
        RECT 794.405 45.940 800.795 46.230 ;
        RECT 793.820 45.360 804.475 45.695 ;
        RECT 793.170 44.775 796.090 45.075 ;
        RECT 799.635 44.760 803.005 45.060 ;
        RECT 791.385 44.025 791.765 44.405 ;
        RECT 793.790 44.040 795.570 44.330 ;
        RECT 797.045 44.130 798.235 44.415 ;
        RECT 801.165 44.010 802.475 44.330 ;
        RECT 792.520 43.425 792.900 43.805 ;
        RECT 796.265 43.465 796.645 43.845 ;
        RECT 798.975 43.455 799.355 43.835 ;
        RECT 800.385 43.300 803.565 43.620 ;
        RECT 790.315 40.710 794.410 40.715 ;
        RECT 805.025 40.710 805.405 46.540 ;
        RECT 813.905 46.490 818.405 46.800 ;
        RECT 905.625 46.400 909.755 46.700 ;
        RECT 809.865 45.940 816.255 46.230 ;
        RECT 821.135 46.190 857.045 46.330 ;
        RECT 821.135 46.060 888.410 46.190 ;
        RECT 856.665 45.920 888.410 46.060 ;
        RECT 809.280 45.360 819.785 45.695 ;
        RECT 844.755 45.495 855.305 45.830 ;
        RECT 892.630 45.800 899.020 46.090 ;
        RECT 808.630 44.775 811.550 45.075 ;
        RECT 815.095 44.760 818.465 45.060 ;
        RECT 823.345 44.855 824.650 45.235 ;
        RECT 825.350 44.855 828.650 45.235 ;
        RECT 829.350 44.855 832.650 45.235 ;
        RECT 833.350 44.855 834.710 45.235 ;
        RECT 836.685 44.855 838.150 45.235 ;
        RECT 838.850 44.855 842.150 45.235 ;
        RECT 842.850 44.855 846.150 45.235 ;
        RECT 846.850 44.855 848.030 45.235 ;
        RECT 892.045 45.220 902.525 45.555 ;
        RECT 862.015 44.715 863.320 45.095 ;
        RECT 868.020 44.715 871.320 45.095 ;
        RECT 872.020 44.715 873.380 45.095 ;
        RECT 875.355 44.715 876.820 45.095 ;
        RECT 877.520 44.715 880.820 45.095 ;
        RECT 885.520 44.715 886.700 45.095 ;
        RECT 824.810 44.510 825.190 44.545 ;
        RECT 806.845 44.025 807.225 44.405 ;
        RECT 809.250 44.040 811.030 44.330 ;
        RECT 812.505 44.130 813.695 44.415 ;
        RECT 816.625 44.010 817.935 44.330 ;
        RECT 824.545 44.200 827.555 44.510 ;
        RECT 824.810 44.165 825.190 44.200 ;
        RECT 828.810 44.165 829.900 44.545 ;
        RECT 832.810 44.540 833.190 44.545 ;
        RECT 830.330 44.175 833.195 44.540 ;
        RECT 838.310 44.520 838.690 44.545 ;
        RECT 838.295 44.200 840.440 44.520 ;
        RECT 832.810 44.165 833.190 44.175 ;
        RECT 838.310 44.165 838.690 44.200 ;
        RECT 841.355 44.165 842.690 44.545 ;
        RECT 846.310 44.525 846.690 44.545 ;
        RECT 843.845 44.205 846.755 44.525 ;
        RECT 863.480 44.370 863.860 44.405 ;
        RECT 846.310 44.165 846.690 44.205 ;
        RECT 863.215 44.060 866.225 44.370 ;
        RECT 863.480 44.025 863.860 44.060 ;
        RECT 867.480 44.025 868.570 44.405 ;
        RECT 871.480 44.400 871.860 44.405 ;
        RECT 869.000 44.035 871.865 44.400 ;
        RECT 876.980 44.380 877.360 44.405 ;
        RECT 876.965 44.060 879.110 44.380 ;
        RECT 871.480 44.025 871.860 44.035 ;
        RECT 876.980 44.025 877.360 44.060 ;
        RECT 880.025 44.025 881.360 44.405 ;
        RECT 884.980 44.385 885.360 44.405 ;
        RECT 882.515 44.065 885.425 44.385 ;
        RECT 884.980 44.025 885.360 44.065 ;
        RECT 889.610 43.885 889.990 44.265 ;
        RECT 892.015 43.900 893.795 44.190 ;
        RECT 895.270 43.990 896.460 44.275 ;
        RECT 899.390 43.870 900.700 44.190 ;
        RECT 807.980 43.425 808.360 43.805 ;
        RECT 811.725 43.465 812.105 43.845 ;
        RECT 814.435 43.455 814.815 43.835 ;
        RECT 815.845 43.300 819.025 43.620 ;
        RECT 890.745 43.285 891.125 43.665 ;
        RECT 894.490 43.325 894.870 43.705 ;
        RECT 897.200 43.315 897.580 43.695 ;
        RECT 823.160 42.855 824.650 43.235 ;
        RECT 825.350 42.855 826.635 43.235 ;
        RECT 844.665 42.855 846.150 43.235 ;
        RECT 846.850 42.855 847.925 43.235 ;
        RECT 898.610 43.160 901.790 43.480 ;
        RECT 861.830 42.715 863.320 43.095 ;
        RECT 885.520 42.715 886.595 43.095 ;
        RECT 824.810 42.165 825.900 42.545 ;
        RECT 826.855 42.175 828.375 42.535 ;
        RECT 829.295 42.170 842.145 42.505 ;
        RECT 846.310 42.500 846.690 42.545 ;
        RECT 845.575 42.200 846.885 42.500 ;
        RECT 846.310 42.165 846.690 42.200 ;
        RECT 863.480 42.025 864.570 42.405 ;
        RECT 865.525 42.035 867.045 42.395 ;
        RECT 867.965 42.030 880.815 42.365 ;
        RECT 884.980 42.360 885.360 42.405 ;
        RECT 884.245 42.060 885.555 42.360 ;
        RECT 884.980 42.025 885.360 42.060 ;
        RECT 821.665 41.530 854.745 41.655 ;
        RECT 821.665 41.305 886.990 41.530 ;
        RECT 854.040 41.165 886.990 41.305 ;
        RECT 888.785 41.155 893.045 41.510 ;
        RECT 805.775 40.710 809.870 40.715 ;
        RECT 789.195 40.705 794.410 40.710 ;
        RECT 804.655 40.705 809.870 40.710 ;
        RECT 820.115 40.705 860.365 40.710 ;
        RECT 789.195 40.570 860.365 40.705 ;
        RECT 886.990 40.570 892.635 40.575 ;
        RECT 903.250 40.570 903.630 46.400 ;
        RECT 912.130 46.350 916.630 46.660 ;
        RECT 988.280 46.540 992.410 46.840 ;
        RECT 908.090 45.800 914.480 46.090 ;
        RECT 907.505 45.220 923.525 45.555 ;
        RECT 972.290 45.495 978.205 45.830 ;
        RECT 975.560 45.475 978.205 45.495 ;
        RECT 906.855 44.635 909.775 44.935 ;
        RECT 913.320 44.620 916.690 44.920 ;
        RECT 952.885 44.855 956.185 45.235 ;
        RECT 956.885 44.855 960.185 45.235 ;
        RECT 966.385 44.855 969.685 45.235 ;
        RECT 970.385 44.855 973.685 45.235 ;
        RECT 905.070 43.885 905.450 44.265 ;
        RECT 907.475 43.900 909.255 44.190 ;
        RECT 910.730 43.990 911.920 44.275 ;
        RECT 914.850 43.870 916.160 44.190 ;
        RECT 906.205 43.285 906.585 43.665 ;
        RECT 909.950 43.325 910.330 43.705 ;
        RECT 912.660 43.315 913.040 43.695 ;
        RECT 914.070 43.160 917.250 43.480 ;
        RECT 952.885 42.855 954.170 43.235 ;
        RECT 972.200 42.855 973.685 43.235 ;
        RECT 904.350 42.075 908.500 42.345 ;
        RECT 954.390 42.175 955.910 42.535 ;
        RECT 985.905 40.710 986.285 46.540 ;
        RECT 994.785 46.490 999.285 46.800 ;
        RECT 1003.740 46.540 1007.870 46.840 ;
        RECT 990.745 45.940 997.135 46.230 ;
        RECT 990.160 45.360 1000.815 45.695 ;
        RECT 989.510 44.775 992.430 45.075 ;
        RECT 995.975 44.760 999.345 45.060 ;
        RECT 987.725 44.025 988.105 44.405 ;
        RECT 990.130 44.040 991.910 44.330 ;
        RECT 993.385 44.130 994.575 44.415 ;
        RECT 997.505 44.010 998.815 44.330 ;
        RECT 988.860 43.425 989.240 43.805 ;
        RECT 992.605 43.465 992.985 43.845 ;
        RECT 995.315 43.455 995.695 43.835 ;
        RECT 996.725 43.300 999.905 43.620 ;
        RECT 986.655 40.710 990.750 40.715 ;
        RECT 1001.365 40.710 1001.745 46.540 ;
        RECT 1010.245 46.490 1014.745 46.800 ;
        RECT 1101.965 46.400 1106.095 46.700 ;
        RECT 1006.205 45.940 1012.595 46.230 ;
        RECT 1017.475 46.190 1053.385 46.330 ;
        RECT 1017.475 46.060 1084.750 46.190 ;
        RECT 1053.005 45.920 1084.750 46.060 ;
        RECT 1005.620 45.360 1016.125 45.695 ;
        RECT 1041.095 45.495 1051.645 45.830 ;
        RECT 1088.970 45.800 1095.360 46.090 ;
        RECT 1004.970 44.775 1007.890 45.075 ;
        RECT 1011.435 44.760 1014.805 45.060 ;
        RECT 1019.685 44.855 1020.990 45.235 ;
        RECT 1021.690 44.855 1024.990 45.235 ;
        RECT 1025.690 44.855 1028.990 45.235 ;
        RECT 1029.690 44.855 1031.050 45.235 ;
        RECT 1033.025 44.855 1034.490 45.235 ;
        RECT 1035.190 44.855 1038.490 45.235 ;
        RECT 1039.190 44.855 1042.490 45.235 ;
        RECT 1043.190 44.855 1044.370 45.235 ;
        RECT 1088.385 45.220 1098.865 45.555 ;
        RECT 1058.355 44.715 1059.660 45.095 ;
        RECT 1064.360 44.715 1067.660 45.095 ;
        RECT 1068.360 44.715 1069.720 45.095 ;
        RECT 1071.695 44.715 1073.160 45.095 ;
        RECT 1073.860 44.715 1077.160 45.095 ;
        RECT 1081.860 44.715 1083.040 45.095 ;
        RECT 1021.150 44.510 1021.530 44.545 ;
        RECT 1003.185 44.025 1003.565 44.405 ;
        RECT 1005.590 44.040 1007.370 44.330 ;
        RECT 1008.845 44.130 1010.035 44.415 ;
        RECT 1012.965 44.010 1014.275 44.330 ;
        RECT 1020.885 44.200 1023.895 44.510 ;
        RECT 1021.150 44.165 1021.530 44.200 ;
        RECT 1025.150 44.165 1026.240 44.545 ;
        RECT 1029.150 44.540 1029.530 44.545 ;
        RECT 1026.670 44.175 1029.535 44.540 ;
        RECT 1034.650 44.520 1035.030 44.545 ;
        RECT 1034.635 44.200 1036.780 44.520 ;
        RECT 1029.150 44.165 1029.530 44.175 ;
        RECT 1034.650 44.165 1035.030 44.200 ;
        RECT 1037.695 44.165 1039.030 44.545 ;
        RECT 1042.650 44.525 1043.030 44.545 ;
        RECT 1040.185 44.205 1043.095 44.525 ;
        RECT 1059.820 44.370 1060.200 44.405 ;
        RECT 1042.650 44.165 1043.030 44.205 ;
        RECT 1059.555 44.060 1062.565 44.370 ;
        RECT 1059.820 44.025 1060.200 44.060 ;
        RECT 1063.820 44.025 1064.910 44.405 ;
        RECT 1067.820 44.400 1068.200 44.405 ;
        RECT 1065.340 44.035 1068.205 44.400 ;
        RECT 1073.320 44.380 1073.700 44.405 ;
        RECT 1073.305 44.060 1075.450 44.380 ;
        RECT 1067.820 44.025 1068.200 44.035 ;
        RECT 1073.320 44.025 1073.700 44.060 ;
        RECT 1076.365 44.025 1077.700 44.405 ;
        RECT 1081.320 44.385 1081.700 44.405 ;
        RECT 1078.855 44.065 1081.765 44.385 ;
        RECT 1081.320 44.025 1081.700 44.065 ;
        RECT 1085.950 43.885 1086.330 44.265 ;
        RECT 1088.355 43.900 1090.135 44.190 ;
        RECT 1091.610 43.990 1092.800 44.275 ;
        RECT 1095.730 43.870 1097.040 44.190 ;
        RECT 1004.320 43.425 1004.700 43.805 ;
        RECT 1008.065 43.465 1008.445 43.845 ;
        RECT 1010.775 43.455 1011.155 43.835 ;
        RECT 1012.185 43.300 1015.365 43.620 ;
        RECT 1087.085 43.285 1087.465 43.665 ;
        RECT 1090.830 43.325 1091.210 43.705 ;
        RECT 1093.540 43.315 1093.920 43.695 ;
        RECT 1019.500 42.855 1020.990 43.235 ;
        RECT 1021.690 42.855 1022.975 43.235 ;
        RECT 1041.005 42.855 1042.490 43.235 ;
        RECT 1043.190 42.855 1044.265 43.235 ;
        RECT 1094.950 43.160 1098.130 43.480 ;
        RECT 1058.170 42.715 1059.660 43.095 ;
        RECT 1081.860 42.715 1082.935 43.095 ;
        RECT 1021.150 42.165 1022.240 42.545 ;
        RECT 1023.195 42.175 1024.715 42.535 ;
        RECT 1025.635 42.170 1038.485 42.505 ;
        RECT 1042.650 42.500 1043.030 42.545 ;
        RECT 1041.915 42.200 1043.225 42.500 ;
        RECT 1042.650 42.165 1043.030 42.200 ;
        RECT 1059.820 42.025 1060.910 42.405 ;
        RECT 1061.865 42.035 1063.385 42.395 ;
        RECT 1064.305 42.030 1077.155 42.365 ;
        RECT 1081.320 42.360 1081.700 42.405 ;
        RECT 1080.585 42.060 1081.895 42.360 ;
        RECT 1081.320 42.025 1081.700 42.060 ;
        RECT 1018.005 41.530 1051.085 41.655 ;
        RECT 1018.005 41.305 1083.330 41.530 ;
        RECT 1050.380 41.165 1083.330 41.305 ;
        RECT 1085.125 41.155 1089.385 41.510 ;
        RECT 1002.115 40.710 1006.210 40.715 ;
        RECT 904.000 40.570 908.095 40.575 ;
        RECT 789.195 40.565 892.635 40.570 ;
        RECT 902.880 40.565 908.095 40.570 ;
        RECT 789.195 39.810 917.910 40.565 ;
        RECT 949.200 39.810 975.855 40.710 ;
        RECT 985.535 40.705 990.750 40.710 ;
        RECT 1000.995 40.705 1006.210 40.710 ;
        RECT 1016.455 40.705 1056.705 40.710 ;
        RECT 985.535 40.570 1056.705 40.705 ;
        RECT 1083.330 40.570 1088.975 40.575 ;
        RECT 1099.590 40.570 1099.970 46.400 ;
        RECT 1108.470 46.350 1112.970 46.660 ;
        RECT 1184.620 46.540 1188.750 46.840 ;
        RECT 1104.430 45.800 1110.820 46.090 ;
        RECT 1103.845 45.220 1119.865 45.555 ;
        RECT 1168.615 45.500 1174.530 45.835 ;
        RECT 1171.885 45.480 1174.530 45.500 ;
        RECT 1103.195 44.635 1106.115 44.935 ;
        RECT 1109.660 44.620 1113.030 44.920 ;
        RECT 1149.210 44.860 1152.510 45.240 ;
        RECT 1153.210 44.860 1156.510 45.240 ;
        RECT 1162.710 44.860 1166.010 45.240 ;
        RECT 1166.710 44.860 1170.010 45.240 ;
        RECT 1101.410 43.885 1101.790 44.265 ;
        RECT 1103.815 43.900 1105.595 44.190 ;
        RECT 1107.070 43.990 1108.260 44.275 ;
        RECT 1111.190 43.870 1112.500 44.190 ;
        RECT 1102.545 43.285 1102.925 43.665 ;
        RECT 1106.290 43.325 1106.670 43.705 ;
        RECT 1109.000 43.315 1109.380 43.695 ;
        RECT 1110.410 43.160 1113.590 43.480 ;
        RECT 1149.210 42.860 1150.495 43.240 ;
        RECT 1168.525 42.860 1170.010 43.240 ;
        RECT 1100.690 42.075 1104.840 42.345 ;
        RECT 1150.715 42.180 1152.235 42.540 ;
        RECT 1100.340 40.570 1104.435 40.575 ;
        RECT 985.535 40.565 1088.975 40.570 ;
        RECT 1099.220 40.565 1104.435 40.570 ;
        RECT 985.535 39.810 1114.250 40.565 ;
        RECT 1145.525 39.815 1172.180 40.715 ;
        RECT 1182.245 40.710 1182.625 46.540 ;
        RECT 1191.125 46.490 1195.625 46.800 ;
        RECT 1200.080 46.540 1204.210 46.840 ;
        RECT 1187.085 45.940 1193.475 46.230 ;
        RECT 1186.500 45.360 1197.155 45.695 ;
        RECT 1185.850 44.775 1188.770 45.075 ;
        RECT 1192.315 44.760 1195.685 45.060 ;
        RECT 1184.065 44.025 1184.445 44.405 ;
        RECT 1186.470 44.040 1188.250 44.330 ;
        RECT 1189.725 44.130 1190.915 44.415 ;
        RECT 1193.845 44.010 1195.155 44.330 ;
        RECT 1185.200 43.425 1185.580 43.805 ;
        RECT 1188.945 43.465 1189.325 43.845 ;
        RECT 1191.655 43.455 1192.035 43.835 ;
        RECT 1193.065 43.300 1196.245 43.620 ;
        RECT 1182.995 40.710 1187.090 40.715 ;
        RECT 1197.705 40.710 1198.085 46.540 ;
        RECT 1206.585 46.490 1211.085 46.800 ;
        RECT 1282.845 46.400 1286.975 46.700 ;
        RECT 1289.350 46.350 1293.850 46.660 ;
        RECT 1298.305 46.400 1302.435 46.700 ;
        RECT 1202.545 45.940 1208.935 46.230 ;
        RECT 1213.815 46.190 1249.725 46.330 ;
        RECT 1213.815 46.060 1281.090 46.190 ;
        RECT 1249.345 45.920 1281.090 46.060 ;
        RECT 1201.960 45.360 1212.465 45.695 ;
        RECT 1237.435 45.495 1247.985 45.830 ;
        RECT 1285.310 45.800 1291.700 46.090 ;
        RECT 1276.105 45.355 1280.050 45.690 ;
        RECT 1201.310 44.775 1204.230 45.075 ;
        RECT 1207.775 44.760 1211.145 45.060 ;
        RECT 1216.025 44.855 1217.330 45.235 ;
        RECT 1218.030 44.855 1221.330 45.235 ;
        RECT 1222.030 44.855 1225.330 45.235 ;
        RECT 1226.030 44.855 1227.390 45.235 ;
        RECT 1229.365 44.855 1230.830 45.235 ;
        RECT 1231.530 44.855 1234.830 45.235 ;
        RECT 1235.530 44.855 1238.830 45.235 ;
        RECT 1239.530 44.855 1240.710 45.235 ;
        RECT 1284.725 45.220 1295.205 45.555 ;
        RECT 1254.695 44.715 1256.000 45.095 ;
        RECT 1256.700 44.715 1260.000 45.095 ;
        RECT 1260.700 44.715 1264.000 45.095 ;
        RECT 1264.700 44.715 1266.060 45.095 ;
        RECT 1268.035 44.715 1269.500 45.095 ;
        RECT 1270.200 44.715 1273.500 45.095 ;
        RECT 1274.200 44.715 1277.500 45.095 ;
        RECT 1278.200 44.715 1279.380 45.095 ;
        RECT 1284.075 44.635 1286.995 44.935 ;
        RECT 1290.540 44.620 1293.910 44.920 ;
        RECT 1217.490 44.510 1217.870 44.545 ;
        RECT 1199.525 44.025 1199.905 44.405 ;
        RECT 1201.930 44.040 1203.710 44.330 ;
        RECT 1205.185 44.130 1206.375 44.415 ;
        RECT 1209.305 44.010 1210.615 44.330 ;
        RECT 1217.225 44.200 1220.235 44.510 ;
        RECT 1217.490 44.165 1217.870 44.200 ;
        RECT 1221.490 44.165 1222.580 44.545 ;
        RECT 1225.490 44.540 1225.870 44.545 ;
        RECT 1223.010 44.175 1225.875 44.540 ;
        RECT 1230.990 44.520 1231.370 44.545 ;
        RECT 1230.975 44.200 1233.120 44.520 ;
        RECT 1225.490 44.165 1225.870 44.175 ;
        RECT 1230.990 44.165 1231.370 44.200 ;
        RECT 1234.035 44.165 1235.370 44.545 ;
        RECT 1238.990 44.525 1239.370 44.545 ;
        RECT 1236.525 44.205 1239.435 44.525 ;
        RECT 1256.160 44.370 1256.540 44.405 ;
        RECT 1238.990 44.165 1239.370 44.205 ;
        RECT 1255.895 44.060 1258.905 44.370 ;
        RECT 1256.160 44.025 1256.540 44.060 ;
        RECT 1260.160 44.025 1261.250 44.405 ;
        RECT 1264.160 44.400 1264.540 44.405 ;
        RECT 1261.680 44.035 1264.545 44.400 ;
        RECT 1269.660 44.380 1270.040 44.405 ;
        RECT 1269.645 44.060 1271.790 44.380 ;
        RECT 1264.160 44.025 1264.540 44.035 ;
        RECT 1269.660 44.025 1270.040 44.060 ;
        RECT 1272.705 44.025 1274.040 44.405 ;
        RECT 1277.660 44.385 1278.040 44.405 ;
        RECT 1275.195 44.065 1278.105 44.385 ;
        RECT 1277.660 44.025 1278.040 44.065 ;
        RECT 1282.290 43.885 1282.670 44.265 ;
        RECT 1284.695 43.900 1286.475 44.190 ;
        RECT 1287.950 43.990 1289.140 44.275 ;
        RECT 1292.070 43.870 1293.380 44.190 ;
        RECT 1200.660 43.425 1201.040 43.805 ;
        RECT 1204.405 43.465 1204.785 43.845 ;
        RECT 1207.115 43.455 1207.495 43.835 ;
        RECT 1208.525 43.300 1211.705 43.620 ;
        RECT 1283.425 43.285 1283.805 43.665 ;
        RECT 1287.170 43.325 1287.550 43.705 ;
        RECT 1289.880 43.315 1290.260 43.695 ;
        RECT 1215.840 42.855 1217.330 43.235 ;
        RECT 1218.030 42.855 1219.315 43.235 ;
        RECT 1237.345 42.855 1238.830 43.235 ;
        RECT 1239.530 42.855 1240.605 43.235 ;
        RECT 1291.290 43.160 1294.470 43.480 ;
        RECT 1254.510 42.715 1256.000 43.095 ;
        RECT 1256.700 42.715 1257.985 43.095 ;
        RECT 1276.015 42.715 1277.500 43.095 ;
        RECT 1278.200 42.715 1279.275 43.095 ;
        RECT 1217.490 42.165 1218.580 42.545 ;
        RECT 1219.535 42.175 1221.055 42.535 ;
        RECT 1221.975 42.170 1234.825 42.505 ;
        RECT 1238.990 42.500 1239.370 42.545 ;
        RECT 1238.255 42.200 1239.565 42.500 ;
        RECT 1238.990 42.165 1239.370 42.200 ;
        RECT 1256.160 42.025 1257.250 42.405 ;
        RECT 1258.205 42.035 1259.725 42.395 ;
        RECT 1260.645 42.030 1273.495 42.365 ;
        RECT 1277.660 42.360 1278.040 42.405 ;
        RECT 1276.925 42.060 1278.235 42.360 ;
        RECT 1277.660 42.025 1278.040 42.060 ;
        RECT 1214.345 41.530 1247.425 41.655 ;
        RECT 1214.345 41.305 1279.670 41.530 ;
        RECT 1246.720 41.165 1279.670 41.305 ;
        RECT 1281.465 41.155 1285.725 41.510 ;
        RECT 1198.455 40.710 1202.550 40.715 ;
        RECT 1181.875 40.705 1187.090 40.710 ;
        RECT 1197.335 40.705 1202.550 40.710 ;
        RECT 1212.795 40.705 1253.045 40.710 ;
        RECT 1181.875 40.570 1253.045 40.705 ;
        RECT 1279.670 40.570 1285.315 40.575 ;
        RECT 1295.930 40.570 1296.310 46.400 ;
        RECT 1304.810 46.350 1309.310 46.660 ;
        RECT 1300.770 45.800 1307.160 46.090 ;
        RECT 1299.535 44.635 1302.455 44.935 ;
        RECT 1306.000 44.620 1309.370 44.920 ;
        RECT 1297.750 43.885 1298.130 44.265 ;
        RECT 1303.410 43.990 1304.600 44.275 ;
        RECT 1302.630 43.325 1303.010 43.705 ;
        RECT 1306.750 43.160 1309.930 43.480 ;
        RECT 1297.030 42.075 1301.180 42.345 ;
        RECT 1296.680 40.570 1300.775 40.575 ;
        RECT 1181.875 40.565 1285.315 40.570 ;
        RECT 1295.560 40.565 1300.775 40.570 ;
        RECT 1181.875 39.810 1310.590 40.565 ;
        RECT 467.620 39.635 525.195 39.775 ;
        RECT 663.995 39.670 721.570 39.810 ;
        RECT 860.335 39.670 917.910 39.810 ;
        RECT 1056.675 39.670 1114.250 39.810 ;
        RECT 1253.015 39.670 1310.590 39.810 ;
        RECT 3.685 35.945 76.075 35.955 ;
        RECT -81.530 34.940 -56.095 35.840 ;
        RECT 3.685 35.055 132.430 35.945 ;
        RECT 164.935 35.110 190.370 36.010 ;
        RECT 200.050 35.945 272.440 35.955 ;
        RECT 200.050 35.055 328.795 35.945 ;
        RECT 361.325 35.070 386.760 35.970 ;
        RECT 396.450 35.895 468.840 35.905 ;
        RECT -79.045 32.760 -77.845 33.140 ;
        RECT -76.090 32.545 -73.815 33.055 ;
        RECT -71.190 32.545 -68.890 33.055 ;
        RECT -66.595 32.545 -64.315 33.055 ;
        RECT -59.520 32.860 -58.285 33.240 ;
        RECT -79.045 30.460 -75.785 30.840 ;
        RECT -75.045 30.460 -71.785 30.840 ;
        RECT -65.545 30.460 -62.285 30.840 ;
        RECT -61.545 30.460 -58.285 30.840 ;
        RECT -78.380 28.875 -56.095 28.885 ;
        RECT -78.380 28.545 -54.555 28.875 ;
        RECT -56.315 28.525 -54.555 28.545 ;
        RECT 4.055 27.895 4.435 35.055 ;
        RECT 5.885 30.840 9.260 31.240 ;
        RECT 9.630 30.600 10.010 30.980 ;
        RECT 12.345 30.640 12.725 31.020 ;
        RECT 16.530 30.590 16.910 30.970 ;
        RECT 6.955 30.175 8.695 30.465 ;
        RECT 10.745 30.125 11.945 30.415 ;
        RECT 13.455 30.095 16.065 30.520 ;
        RECT 17.665 30.190 18.045 30.570 ;
        RECT 5.215 27.955 11.940 28.255 ;
        RECT 15.640 27.655 18.745 27.930 ;
        RECT 19.515 27.895 19.895 35.055 ;
        RECT 76.075 35.045 132.430 35.055 ;
        RECT 36.155 34.060 73.705 34.070 ;
        RECT 36.155 33.785 101.835 34.060 ;
        RECT 73.060 33.775 101.835 33.785 ;
        RECT 103.505 33.755 110.210 34.055 ;
        RECT 39.860 32.875 41.060 33.255 ;
        RECT 42.815 32.660 45.090 33.170 ;
        RECT 47.715 32.660 50.015 33.170 ;
        RECT 52.310 32.660 54.590 33.170 ;
        RECT 59.385 32.975 60.620 33.355 ;
        RECT 76.365 32.865 77.820 33.245 ;
        RECT 60.800 32.620 61.180 32.655 ;
        RECT 81.515 32.650 83.790 33.160 ;
        RECT 86.415 32.650 88.715 33.160 ;
        RECT 91.010 32.650 93.290 33.160 ;
        RECT 100.060 32.965 101.340 33.345 ;
        RECT 39.300 32.515 39.680 32.555 ;
        RECT 39.230 32.210 42.065 32.515 ;
        RECT 58.045 32.310 61.180 32.620 ;
        RECT 99.500 32.610 99.880 32.645 ;
        RECT 78.000 32.505 78.380 32.545 ;
        RECT 60.800 32.275 61.180 32.310 ;
        RECT 39.300 32.175 39.680 32.210 ;
        RECT 77.930 32.200 80.765 32.505 ;
        RECT 96.745 32.300 99.880 32.610 ;
        RECT 99.500 32.265 99.880 32.300 ;
        RECT 78.000 32.165 78.380 32.200 ;
        RECT 21.345 30.800 24.750 31.240 ;
        RECT 25.090 30.600 25.470 30.980 ;
        RECT 27.805 30.640 28.185 31.020 ;
        RECT 31.990 30.590 32.370 30.970 ;
        RECT 39.860 30.575 43.120 30.955 ;
        RECT 43.860 30.575 47.120 30.955 ;
        RECT 53.360 30.575 56.620 30.955 ;
        RECT 57.360 30.575 60.620 30.955 ;
        RECT 22.415 30.175 24.155 30.465 ;
        RECT 26.205 30.125 27.405 30.415 ;
        RECT 28.915 30.095 31.510 30.470 ;
        RECT 33.125 30.190 33.505 30.570 ;
        RECT 76.525 30.565 77.820 30.945 ;
        RECT 82.560 30.565 85.820 30.945 ;
        RECT 86.560 30.565 87.745 30.945 ;
        RECT 90.010 30.565 91.320 30.945 ;
        RECT 92.060 30.565 95.320 30.945 ;
        RECT 100.060 30.565 101.075 30.945 ;
        RECT 104.140 30.810 107.555 31.230 ;
        RECT 107.885 30.590 108.265 30.970 ;
        RECT 110.600 30.630 110.980 31.010 ;
        RECT 114.785 30.580 115.165 30.960 ;
        RECT 39.300 29.875 39.680 30.255 ;
        RECT 43.300 29.875 43.680 30.255 ;
        RECT 47.300 30.210 47.680 30.255 ;
        RECT 52.800 30.210 53.180 30.255 ;
        RECT 47.250 29.895 53.185 30.210 ;
        RECT 47.300 29.875 47.680 29.895 ;
        RECT 52.800 29.875 53.180 29.895 ;
        RECT 56.800 29.875 57.180 30.255 ;
        RECT 60.800 29.875 61.180 30.255 ;
        RECT 78.000 29.865 78.380 30.245 ;
        RECT 82.000 29.865 82.380 30.245 ;
        RECT 86.000 30.200 86.380 30.245 ;
        RECT 91.500 30.200 91.880 30.245 ;
        RECT 85.950 29.885 91.885 30.200 ;
        RECT 86.000 29.865 86.380 29.885 ;
        RECT 91.500 29.865 91.880 29.885 ;
        RECT 95.500 29.865 95.880 30.245 ;
        RECT 99.500 29.865 99.880 30.245 ;
        RECT 105.210 30.165 106.950 30.455 ;
        RECT 109.000 30.115 110.200 30.405 ;
        RECT 111.710 30.075 114.340 30.530 ;
        RECT 115.920 30.180 116.300 30.560 ;
        RECT 70.090 29.240 90.865 29.615 ;
        RECT 40.525 28.660 67.835 29.000 ;
        RECT 20.140 27.955 27.400 28.255 ;
        RECT 5.195 27.335 9.320 27.605 ;
        RECT 20.695 27.420 24.780 27.690 ;
        RECT 31.100 27.655 34.850 27.930 ;
        RECT 69.120 27.885 101.085 28.275 ;
        RECT 113.895 27.645 117.025 27.920 ;
        RECT 117.770 27.885 118.150 35.045 ;
        RECT 167.420 32.930 168.620 33.310 ;
        RECT 119.010 32.585 125.750 32.885 ;
        RECT 170.375 32.715 172.650 33.225 ;
        RECT 175.275 32.715 177.575 33.225 ;
        RECT 179.870 32.715 182.150 33.225 ;
        RECT 186.945 33.030 188.180 33.410 ;
        RECT 119.600 30.790 123.055 31.230 ;
        RECT 123.345 30.590 123.725 30.970 ;
        RECT 126.060 30.630 126.440 31.010 ;
        RECT 130.245 30.580 130.625 30.960 ;
        RECT 167.420 30.630 170.680 31.010 ;
        RECT 171.420 30.630 174.680 31.010 ;
        RECT 180.920 30.630 184.180 31.010 ;
        RECT 184.920 30.630 188.180 31.010 ;
        RECT 120.670 30.165 122.410 30.455 ;
        RECT 124.460 30.115 125.660 30.405 ;
        RECT 127.170 30.085 129.795 30.495 ;
        RECT 131.380 30.180 131.760 30.560 ;
        RECT 118.415 29.405 134.335 29.705 ;
        RECT 168.085 28.980 190.370 29.055 ;
        RECT 118.950 28.660 135.895 28.960 ;
        RECT 168.085 28.715 194.430 28.980 ;
        RECT 190.255 28.640 194.430 28.715 ;
        RECT 129.355 27.645 137.055 27.920 ;
        RECT 200.420 27.895 200.800 35.055 ;
        RECT 202.250 30.840 205.625 31.240 ;
        RECT 205.995 30.600 206.375 30.980 ;
        RECT 208.710 30.640 209.090 31.020 ;
        RECT 212.895 30.590 213.275 30.970 ;
        RECT 203.320 30.175 205.060 30.465 ;
        RECT 207.110 30.125 208.310 30.415 ;
        RECT 209.820 30.095 212.430 30.520 ;
        RECT 214.030 30.190 214.410 30.570 ;
        RECT 201.565 29.415 215.130 29.730 ;
        RECT 201.560 28.670 215.120 28.970 ;
        RECT 201.580 27.955 208.305 28.255 ;
        RECT 212.005 27.655 215.110 27.930 ;
        RECT 215.880 27.895 216.260 35.055 ;
        RECT 272.440 35.045 328.795 35.055 ;
        RECT 232.520 34.060 270.070 34.070 ;
        RECT 232.520 33.785 298.200 34.060 ;
        RECT 269.425 33.775 298.200 33.785 ;
        RECT 299.870 33.755 306.575 34.055 ;
        RECT 234.030 32.875 235.485 33.255 ;
        RECT 236.225 32.875 237.425 33.255 ;
        RECT 239.180 32.660 241.455 33.170 ;
        RECT 244.080 32.660 246.380 33.170 ;
        RECT 248.675 32.660 250.955 33.170 ;
        RECT 255.750 32.975 256.985 33.355 ;
        RECT 257.725 32.975 259.005 33.355 ;
        RECT 272.730 32.865 274.185 33.245 ;
        RECT 257.165 32.620 257.545 32.655 ;
        RECT 277.880 32.650 280.155 33.160 ;
        RECT 282.780 32.650 285.080 33.160 ;
        RECT 287.375 32.650 289.655 33.160 ;
        RECT 296.425 32.965 297.705 33.345 ;
        RECT 235.665 32.515 236.045 32.555 ;
        RECT 235.595 32.210 238.430 32.515 ;
        RECT 254.410 32.310 257.545 32.620 ;
        RECT 295.865 32.610 296.245 32.645 ;
        RECT 274.365 32.505 274.745 32.545 ;
        RECT 257.165 32.275 257.545 32.310 ;
        RECT 235.665 32.175 236.045 32.210 ;
        RECT 274.295 32.200 277.130 32.505 ;
        RECT 293.110 32.300 296.245 32.610 ;
        RECT 295.865 32.265 296.245 32.300 ;
        RECT 274.365 32.165 274.745 32.200 ;
        RECT 217.710 30.800 221.115 31.240 ;
        RECT 221.455 30.600 221.835 30.980 ;
        RECT 224.170 30.640 224.550 31.020 ;
        RECT 228.355 30.590 228.735 30.970 ;
        RECT 234.190 30.575 235.485 30.955 ;
        RECT 236.225 30.575 239.485 30.955 ;
        RECT 240.225 30.575 243.485 30.955 ;
        RECT 244.225 30.575 245.410 30.955 ;
        RECT 247.675 30.575 248.985 30.955 ;
        RECT 249.725 30.575 252.985 30.955 ;
        RECT 253.725 30.575 256.985 30.955 ;
        RECT 257.725 30.575 258.740 30.955 ;
        RECT 218.780 30.175 220.520 30.465 ;
        RECT 222.570 30.125 223.770 30.415 ;
        RECT 225.280 30.095 227.875 30.470 ;
        RECT 229.490 30.190 229.870 30.570 ;
        RECT 272.890 30.565 274.185 30.945 ;
        RECT 278.925 30.565 282.185 30.945 ;
        RECT 282.925 30.565 284.110 30.945 ;
        RECT 286.375 30.565 287.685 30.945 ;
        RECT 288.425 30.565 291.685 30.945 ;
        RECT 296.425 30.565 297.440 30.945 ;
        RECT 300.505 30.810 303.920 31.230 ;
        RECT 304.250 30.590 304.630 30.970 ;
        RECT 306.965 30.630 307.345 31.010 ;
        RECT 311.150 30.580 311.530 30.960 ;
        RECT 235.665 29.875 236.045 30.255 ;
        RECT 239.665 29.875 240.045 30.255 ;
        RECT 243.665 30.210 244.045 30.255 ;
        RECT 249.165 30.210 249.545 30.255 ;
        RECT 243.615 29.895 249.550 30.210 ;
        RECT 243.665 29.875 244.045 29.895 ;
        RECT 249.165 29.875 249.545 29.895 ;
        RECT 253.165 29.875 253.545 30.255 ;
        RECT 257.165 29.875 257.545 30.255 ;
        RECT 274.365 29.865 274.745 30.245 ;
        RECT 278.365 29.865 278.745 30.245 ;
        RECT 282.365 30.200 282.745 30.245 ;
        RECT 287.865 30.200 288.245 30.245 ;
        RECT 282.315 29.885 288.250 30.200 ;
        RECT 282.365 29.865 282.745 29.885 ;
        RECT 287.865 29.865 288.245 29.885 ;
        RECT 291.865 29.865 292.245 30.245 ;
        RECT 295.865 29.865 296.245 30.245 ;
        RECT 301.575 30.165 303.315 30.455 ;
        RECT 305.365 30.115 306.565 30.405 ;
        RECT 308.075 30.075 310.705 30.530 ;
        RECT 312.285 30.180 312.665 30.560 ;
        RECT 217.020 29.415 230.845 29.715 ;
        RECT 232.520 29.250 248.530 29.625 ;
        RECT 266.455 29.240 287.230 29.615 ;
        RECT 217.025 28.670 235.445 28.970 ;
        RECT 236.890 28.660 264.200 29.000 ;
        RECT 216.505 27.955 223.765 28.255 ;
        RECT 36.155 27.530 54.825 27.540 ;
        RECT 36.155 27.520 93.525 27.530 ;
        RECT 36.155 27.220 102.530 27.520 ;
        RECT 201.560 27.335 205.685 27.605 ;
        RECT 217.060 27.420 221.145 27.690 ;
        RECT 227.465 27.655 231.215 27.930 ;
        RECT 232.520 27.895 258.750 28.285 ;
        RECT 265.485 27.885 297.450 28.275 ;
        RECT 310.260 27.645 313.390 27.920 ;
        RECT 314.135 27.885 314.515 35.045 ;
        RECT 396.450 35.005 525.195 35.895 ;
        RECT 557.645 35.115 583.080 36.015 ;
        RECT 592.825 35.930 665.215 35.940 ;
        RECT 592.825 35.040 721.570 35.930 ;
        RECT 754.010 35.120 779.445 36.020 ;
        RECT 789.165 35.930 861.555 35.940 ;
        RECT 789.165 35.040 917.910 35.930 ;
        RECT 950.395 35.105 975.830 36.005 ;
        RECT 985.505 35.930 1057.895 35.940 ;
        RECT 985.505 35.040 1114.250 35.930 ;
        RECT 1146.720 35.110 1172.155 36.010 ;
        RECT 1181.845 35.930 1254.235 35.940 ;
        RECT 1181.845 35.040 1310.590 35.930 ;
        RECT 363.810 32.890 365.010 33.270 ;
        RECT 315.375 32.585 322.115 32.885 ;
        RECT 366.765 32.675 369.040 33.185 ;
        RECT 371.665 32.675 373.965 33.185 ;
        RECT 376.260 32.675 378.540 33.185 ;
        RECT 383.335 32.990 384.570 33.370 ;
        RECT 315.965 30.790 319.420 31.230 ;
        RECT 319.710 30.590 320.090 30.970 ;
        RECT 322.425 30.630 322.805 31.010 ;
        RECT 326.610 30.580 326.990 30.960 ;
        RECT 363.810 30.590 367.070 30.970 ;
        RECT 367.810 30.590 371.070 30.970 ;
        RECT 377.310 30.590 380.570 30.970 ;
        RECT 381.310 30.590 384.570 30.970 ;
        RECT 317.035 30.165 318.775 30.455 ;
        RECT 320.825 30.115 322.025 30.405 ;
        RECT 323.535 30.085 326.160 30.495 ;
        RECT 327.745 30.180 328.125 30.560 ;
        RECT 314.780 29.405 330.700 29.705 ;
        RECT 315.315 28.660 332.260 28.960 ;
        RECT 364.475 28.940 386.760 29.015 ;
        RECT 364.475 28.675 390.820 28.940 ;
        RECT 386.645 28.600 390.820 28.675 ;
        RECT 325.720 27.645 333.420 27.920 ;
        RECT 396.820 27.845 397.200 35.005 ;
        RECT 398.650 30.790 402.025 31.190 ;
        RECT 402.395 30.550 402.775 30.930 ;
        RECT 405.110 30.590 405.490 30.970 ;
        RECT 409.295 30.540 409.675 30.920 ;
        RECT 399.720 30.125 401.460 30.415 ;
        RECT 403.510 30.075 404.710 30.365 ;
        RECT 406.220 30.045 408.830 30.470 ;
        RECT 410.430 30.140 410.810 30.520 ;
        RECT 397.965 29.365 411.530 29.680 ;
        RECT 397.960 28.620 411.520 28.920 ;
        RECT 397.980 27.905 404.705 28.205 ;
        RECT 408.405 27.605 411.510 27.880 ;
        RECT 412.280 27.845 412.660 35.005 ;
        RECT 468.840 34.995 525.195 35.005 ;
        RECT 428.920 34.010 466.470 34.020 ;
        RECT 428.920 33.735 494.600 34.010 ;
        RECT 465.825 33.725 494.600 33.735 ;
        RECT 496.270 33.705 502.975 34.005 ;
        RECT 430.430 32.825 431.885 33.205 ;
        RECT 432.625 32.825 433.825 33.205 ;
        RECT 435.580 32.610 437.855 33.120 ;
        RECT 440.480 32.610 442.780 33.120 ;
        RECT 445.075 32.610 447.355 33.120 ;
        RECT 452.150 32.925 453.385 33.305 ;
        RECT 454.125 32.925 455.405 33.305 ;
        RECT 469.130 32.815 470.585 33.195 ;
        RECT 453.565 32.570 453.945 32.605 ;
        RECT 474.280 32.600 476.555 33.110 ;
        RECT 479.180 32.600 481.480 33.110 ;
        RECT 483.775 32.600 486.055 33.110 ;
        RECT 492.825 32.915 494.105 33.295 ;
        RECT 432.065 32.465 432.445 32.505 ;
        RECT 431.995 32.160 434.830 32.465 ;
        RECT 450.810 32.260 453.945 32.570 ;
        RECT 492.265 32.560 492.645 32.595 ;
        RECT 470.765 32.455 471.145 32.495 ;
        RECT 453.565 32.225 453.945 32.260 ;
        RECT 432.065 32.125 432.445 32.160 ;
        RECT 470.695 32.150 473.530 32.455 ;
        RECT 489.510 32.250 492.645 32.560 ;
        RECT 492.265 32.215 492.645 32.250 ;
        RECT 470.765 32.115 471.145 32.150 ;
        RECT 414.110 30.750 417.515 31.190 ;
        RECT 417.855 30.550 418.235 30.930 ;
        RECT 420.570 30.590 420.950 30.970 ;
        RECT 424.755 30.540 425.135 30.920 ;
        RECT 430.590 30.525 431.885 30.905 ;
        RECT 432.625 30.525 435.885 30.905 ;
        RECT 436.625 30.525 439.885 30.905 ;
        RECT 440.625 30.525 441.810 30.905 ;
        RECT 444.075 30.525 445.385 30.905 ;
        RECT 446.125 30.525 449.385 30.905 ;
        RECT 450.125 30.525 453.385 30.905 ;
        RECT 454.125 30.525 455.140 30.905 ;
        RECT 415.180 30.125 416.920 30.415 ;
        RECT 418.970 30.075 420.170 30.365 ;
        RECT 421.680 30.045 424.275 30.420 ;
        RECT 425.890 30.140 426.270 30.520 ;
        RECT 469.290 30.515 470.585 30.895 ;
        RECT 475.325 30.515 478.585 30.895 ;
        RECT 479.325 30.515 480.510 30.895 ;
        RECT 482.775 30.515 484.085 30.895 ;
        RECT 484.825 30.515 488.085 30.895 ;
        RECT 492.825 30.515 493.840 30.895 ;
        RECT 496.905 30.760 500.320 31.180 ;
        RECT 500.650 30.540 501.030 30.920 ;
        RECT 503.365 30.580 503.745 30.960 ;
        RECT 507.550 30.530 507.930 30.910 ;
        RECT 432.065 29.825 432.445 30.205 ;
        RECT 436.065 29.825 436.445 30.205 ;
        RECT 440.065 30.160 440.445 30.205 ;
        RECT 445.565 30.160 445.945 30.205 ;
        RECT 440.015 29.845 445.950 30.160 ;
        RECT 440.065 29.825 440.445 29.845 ;
        RECT 445.565 29.825 445.945 29.845 ;
        RECT 449.565 29.825 449.945 30.205 ;
        RECT 453.565 29.825 453.945 30.205 ;
        RECT 470.765 29.815 471.145 30.195 ;
        RECT 474.765 29.815 475.145 30.195 ;
        RECT 478.765 30.150 479.145 30.195 ;
        RECT 484.265 30.150 484.645 30.195 ;
        RECT 478.715 29.835 484.650 30.150 ;
        RECT 478.765 29.815 479.145 29.835 ;
        RECT 484.265 29.815 484.645 29.835 ;
        RECT 488.265 29.815 488.645 30.195 ;
        RECT 492.265 29.815 492.645 30.195 ;
        RECT 497.975 30.115 499.715 30.405 ;
        RECT 501.765 30.065 502.965 30.355 ;
        RECT 504.475 30.025 507.105 30.480 ;
        RECT 508.685 30.130 509.065 30.510 ;
        RECT 413.420 29.365 427.245 29.665 ;
        RECT 428.920 29.200 444.930 29.575 ;
        RECT 462.855 29.190 483.630 29.565 ;
        RECT 413.425 28.620 431.845 28.920 ;
        RECT 433.290 28.610 460.600 28.950 ;
        RECT 412.905 27.905 420.165 28.205 ;
        RECT 232.520 27.530 251.190 27.540 ;
        RECT 232.520 27.520 289.890 27.530 ;
        RECT 232.520 27.220 298.895 27.520 ;
        RECT 397.960 27.285 402.085 27.555 ;
        RECT 413.460 27.370 417.545 27.640 ;
        RECT 423.865 27.605 427.615 27.880 ;
        RECT 428.920 27.845 455.150 28.235 ;
        RECT 461.885 27.835 493.850 28.225 ;
        RECT 506.660 27.595 509.790 27.870 ;
        RECT 510.535 27.835 510.915 34.995 ;
        RECT 560.130 32.935 561.330 33.315 ;
        RECT 511.775 32.535 518.515 32.835 ;
        RECT 563.085 32.720 565.360 33.230 ;
        RECT 567.985 32.720 570.285 33.230 ;
        RECT 572.580 32.720 574.860 33.230 ;
        RECT 579.655 33.035 580.890 33.415 ;
        RECT 512.365 30.740 515.820 31.180 ;
        RECT 516.110 30.540 516.490 30.920 ;
        RECT 518.825 30.580 519.205 30.960 ;
        RECT 523.010 30.530 523.390 30.910 ;
        RECT 560.130 30.635 563.390 31.015 ;
        RECT 564.130 30.635 567.390 31.015 ;
        RECT 573.630 30.635 576.890 31.015 ;
        RECT 577.630 30.635 580.890 31.015 ;
        RECT 513.435 30.115 515.175 30.405 ;
        RECT 517.225 30.065 518.425 30.355 ;
        RECT 519.935 30.035 522.560 30.445 ;
        RECT 524.145 30.130 524.525 30.510 ;
        RECT 511.180 29.355 527.100 29.655 ;
        RECT 560.795 28.985 583.080 29.060 ;
        RECT 511.715 28.610 528.660 28.910 ;
        RECT 560.795 28.720 587.140 28.985 ;
        RECT 582.965 28.645 587.140 28.720 ;
        RECT 593.195 27.880 593.575 35.040 ;
        RECT 595.025 30.825 598.400 31.225 ;
        RECT 598.770 30.585 599.150 30.965 ;
        RECT 601.485 30.625 601.865 31.005 ;
        RECT 605.670 30.575 606.050 30.955 ;
        RECT 596.095 30.160 597.835 30.450 ;
        RECT 599.885 30.110 601.085 30.400 ;
        RECT 602.595 30.080 605.205 30.505 ;
        RECT 606.805 30.175 607.185 30.555 ;
        RECT 594.340 29.400 607.905 29.715 ;
        RECT 594.335 28.655 607.895 28.955 ;
        RECT 594.355 27.940 601.080 28.240 ;
        RECT 522.120 27.595 529.820 27.870 ;
        RECT 604.780 27.640 607.885 27.915 ;
        RECT 608.655 27.880 609.035 35.040 ;
        RECT 665.215 35.030 721.570 35.040 ;
        RECT 625.295 34.045 662.845 34.055 ;
        RECT 625.295 33.770 690.975 34.045 ;
        RECT 662.200 33.760 690.975 33.770 ;
        RECT 692.645 33.740 699.350 34.040 ;
        RECT 626.805 32.860 628.260 33.240 ;
        RECT 629.000 32.860 630.200 33.240 ;
        RECT 631.955 32.645 634.230 33.155 ;
        RECT 636.855 32.645 639.155 33.155 ;
        RECT 641.450 32.645 643.730 33.155 ;
        RECT 648.525 32.960 649.760 33.340 ;
        RECT 650.500 32.960 651.780 33.340 ;
        RECT 665.505 32.850 666.960 33.230 ;
        RECT 649.940 32.605 650.320 32.640 ;
        RECT 670.655 32.635 672.930 33.145 ;
        RECT 675.555 32.635 677.855 33.145 ;
        RECT 680.150 32.635 682.430 33.145 ;
        RECT 689.200 32.950 690.480 33.330 ;
        RECT 628.440 32.500 628.820 32.540 ;
        RECT 628.370 32.195 631.205 32.500 ;
        RECT 647.185 32.295 650.320 32.605 ;
        RECT 688.640 32.595 689.020 32.630 ;
        RECT 667.140 32.490 667.520 32.530 ;
        RECT 649.940 32.260 650.320 32.295 ;
        RECT 628.440 32.160 628.820 32.195 ;
        RECT 667.070 32.185 669.905 32.490 ;
        RECT 685.885 32.285 689.020 32.595 ;
        RECT 688.640 32.250 689.020 32.285 ;
        RECT 667.140 32.150 667.520 32.185 ;
        RECT 610.485 30.785 613.890 31.225 ;
        RECT 614.230 30.585 614.610 30.965 ;
        RECT 616.945 30.625 617.325 31.005 ;
        RECT 621.130 30.575 621.510 30.955 ;
        RECT 626.965 30.560 628.260 30.940 ;
        RECT 629.000 30.560 632.260 30.940 ;
        RECT 633.000 30.560 636.260 30.940 ;
        RECT 637.000 30.560 638.185 30.940 ;
        RECT 640.450 30.560 641.760 30.940 ;
        RECT 642.500 30.560 645.760 30.940 ;
        RECT 646.500 30.560 649.760 30.940 ;
        RECT 650.500 30.560 651.515 30.940 ;
        RECT 611.555 30.160 613.295 30.450 ;
        RECT 615.345 30.110 616.545 30.400 ;
        RECT 618.055 30.080 620.650 30.455 ;
        RECT 622.265 30.175 622.645 30.555 ;
        RECT 665.665 30.550 666.960 30.930 ;
        RECT 671.700 30.550 674.960 30.930 ;
        RECT 675.700 30.550 676.885 30.930 ;
        RECT 679.150 30.550 680.460 30.930 ;
        RECT 681.200 30.550 684.460 30.930 ;
        RECT 689.200 30.550 690.215 30.930 ;
        RECT 693.280 30.795 696.695 31.215 ;
        RECT 697.025 30.575 697.405 30.955 ;
        RECT 699.740 30.615 700.120 30.995 ;
        RECT 703.925 30.565 704.305 30.945 ;
        RECT 628.440 29.860 628.820 30.240 ;
        RECT 632.440 29.860 632.820 30.240 ;
        RECT 636.440 30.195 636.820 30.240 ;
        RECT 641.940 30.195 642.320 30.240 ;
        RECT 636.390 29.880 642.325 30.195 ;
        RECT 636.440 29.860 636.820 29.880 ;
        RECT 641.940 29.860 642.320 29.880 ;
        RECT 645.940 29.860 646.320 30.240 ;
        RECT 649.940 29.860 650.320 30.240 ;
        RECT 667.140 29.850 667.520 30.230 ;
        RECT 671.140 29.850 671.520 30.230 ;
        RECT 675.140 30.185 675.520 30.230 ;
        RECT 680.640 30.185 681.020 30.230 ;
        RECT 675.090 29.870 681.025 30.185 ;
        RECT 675.140 29.850 675.520 29.870 ;
        RECT 680.640 29.850 681.020 29.870 ;
        RECT 684.640 29.850 685.020 30.230 ;
        RECT 688.640 29.850 689.020 30.230 ;
        RECT 694.350 30.150 696.090 30.440 ;
        RECT 698.140 30.100 699.340 30.390 ;
        RECT 700.850 30.060 703.480 30.515 ;
        RECT 705.060 30.165 705.440 30.545 ;
        RECT 609.795 29.400 623.620 29.700 ;
        RECT 625.295 29.235 641.305 29.610 ;
        RECT 659.230 29.225 680.005 29.600 ;
        RECT 609.800 28.655 628.220 28.955 ;
        RECT 629.665 28.645 656.975 28.985 ;
        RECT 609.280 27.940 616.540 28.240 ;
        RECT 428.920 27.480 447.590 27.490 ;
        RECT 428.920 27.470 486.290 27.480 ;
        RECT 65.965 27.210 102.530 27.220 ;
        RECT 262.330 27.210 298.895 27.220 ;
        RECT 428.920 27.170 495.295 27.470 ;
        RECT 594.335 27.320 598.460 27.590 ;
        RECT 609.835 27.405 613.920 27.675 ;
        RECT 620.240 27.640 623.990 27.915 ;
        RECT 625.295 27.880 651.525 28.270 ;
        RECT 658.260 27.870 690.225 28.260 ;
        RECT 703.035 27.630 706.165 27.905 ;
        RECT 706.910 27.870 707.290 35.030 ;
        RECT 756.495 32.940 757.695 33.320 ;
        RECT 708.150 32.570 714.890 32.870 ;
        RECT 759.450 32.725 761.725 33.235 ;
        RECT 764.350 32.725 766.650 33.235 ;
        RECT 768.945 32.725 771.225 33.235 ;
        RECT 776.020 33.040 777.255 33.420 ;
        RECT 708.740 30.775 712.195 31.215 ;
        RECT 712.485 30.575 712.865 30.955 ;
        RECT 715.200 30.615 715.580 30.995 ;
        RECT 719.385 30.565 719.765 30.945 ;
        RECT 756.495 30.640 759.755 31.020 ;
        RECT 760.495 30.640 763.755 31.020 ;
        RECT 769.995 30.640 773.255 31.020 ;
        RECT 773.995 30.640 777.255 31.020 ;
        RECT 709.810 30.150 711.550 30.440 ;
        RECT 713.600 30.100 714.800 30.390 ;
        RECT 716.310 30.070 718.935 30.480 ;
        RECT 720.520 30.165 720.900 30.545 ;
        RECT 707.555 29.390 723.475 29.690 ;
        RECT 757.160 28.990 779.445 29.065 ;
        RECT 708.090 28.645 725.035 28.945 ;
        RECT 757.160 28.725 783.505 28.990 ;
        RECT 779.330 28.650 783.505 28.725 ;
        RECT 718.495 27.630 726.195 27.905 ;
        RECT 789.535 27.880 789.915 35.040 ;
        RECT 791.365 30.825 794.740 31.225 ;
        RECT 795.110 30.585 795.490 30.965 ;
        RECT 797.825 30.625 798.205 31.005 ;
        RECT 802.010 30.575 802.390 30.955 ;
        RECT 792.435 30.160 794.175 30.450 ;
        RECT 796.225 30.110 797.425 30.400 ;
        RECT 798.935 30.080 801.545 30.505 ;
        RECT 803.145 30.175 803.525 30.555 ;
        RECT 790.680 29.400 804.245 29.715 ;
        RECT 790.675 28.655 804.235 28.955 ;
        RECT 790.695 27.940 797.420 28.240 ;
        RECT 801.120 27.640 804.225 27.915 ;
        RECT 804.995 27.880 805.375 35.040 ;
        RECT 861.555 35.030 917.910 35.040 ;
        RECT 821.635 34.045 859.185 34.055 ;
        RECT 821.635 33.770 887.315 34.045 ;
        RECT 858.540 33.760 887.315 33.770 ;
        RECT 888.985 33.740 895.690 34.040 ;
        RECT 823.145 32.860 824.600 33.240 ;
        RECT 825.340 32.860 826.540 33.240 ;
        RECT 828.295 32.645 830.570 33.155 ;
        RECT 833.195 32.645 835.495 33.155 ;
        RECT 837.790 32.645 840.070 33.155 ;
        RECT 844.865 32.960 846.100 33.340 ;
        RECT 846.840 32.960 848.120 33.340 ;
        RECT 861.845 32.850 863.300 33.230 ;
        RECT 846.280 32.605 846.660 32.640 ;
        RECT 866.995 32.635 869.270 33.145 ;
        RECT 871.895 32.635 874.195 33.145 ;
        RECT 876.490 32.635 878.770 33.145 ;
        RECT 885.540 32.950 886.820 33.330 ;
        RECT 824.780 32.500 825.160 32.540 ;
        RECT 824.710 32.195 827.545 32.500 ;
        RECT 843.525 32.295 846.660 32.605 ;
        RECT 884.980 32.595 885.360 32.630 ;
        RECT 863.480 32.490 863.860 32.530 ;
        RECT 846.280 32.260 846.660 32.295 ;
        RECT 824.780 32.160 825.160 32.195 ;
        RECT 863.410 32.185 866.245 32.490 ;
        RECT 882.225 32.285 885.360 32.595 ;
        RECT 884.980 32.250 885.360 32.285 ;
        RECT 863.480 32.150 863.860 32.185 ;
        RECT 806.825 30.785 810.230 31.225 ;
        RECT 810.570 30.585 810.950 30.965 ;
        RECT 813.285 30.625 813.665 31.005 ;
        RECT 817.470 30.575 817.850 30.955 ;
        RECT 823.305 30.560 824.600 30.940 ;
        RECT 825.340 30.560 828.600 30.940 ;
        RECT 829.340 30.560 832.600 30.940 ;
        RECT 833.340 30.560 834.525 30.940 ;
        RECT 836.790 30.560 838.100 30.940 ;
        RECT 838.840 30.560 842.100 30.940 ;
        RECT 842.840 30.560 846.100 30.940 ;
        RECT 846.840 30.560 847.855 30.940 ;
        RECT 807.895 30.160 809.635 30.450 ;
        RECT 811.685 30.110 812.885 30.400 ;
        RECT 814.395 30.080 816.990 30.455 ;
        RECT 818.605 30.175 818.985 30.555 ;
        RECT 862.005 30.550 863.300 30.930 ;
        RECT 868.040 30.550 871.300 30.930 ;
        RECT 872.040 30.550 873.225 30.930 ;
        RECT 875.490 30.550 876.800 30.930 ;
        RECT 877.540 30.550 880.800 30.930 ;
        RECT 885.540 30.550 886.555 30.930 ;
        RECT 889.620 30.795 893.035 31.215 ;
        RECT 893.365 30.575 893.745 30.955 ;
        RECT 896.080 30.615 896.460 30.995 ;
        RECT 900.265 30.565 900.645 30.945 ;
        RECT 824.780 29.860 825.160 30.240 ;
        RECT 828.780 29.860 829.160 30.240 ;
        RECT 832.780 30.195 833.160 30.240 ;
        RECT 838.280 30.195 838.660 30.240 ;
        RECT 832.730 29.880 838.665 30.195 ;
        RECT 832.780 29.860 833.160 29.880 ;
        RECT 838.280 29.860 838.660 29.880 ;
        RECT 842.280 29.860 842.660 30.240 ;
        RECT 846.280 29.860 846.660 30.240 ;
        RECT 863.480 29.850 863.860 30.230 ;
        RECT 867.480 29.850 867.860 30.230 ;
        RECT 871.480 30.185 871.860 30.230 ;
        RECT 876.980 30.185 877.360 30.230 ;
        RECT 871.430 29.870 877.365 30.185 ;
        RECT 871.480 29.850 871.860 29.870 ;
        RECT 876.980 29.850 877.360 29.870 ;
        RECT 880.980 29.850 881.360 30.230 ;
        RECT 884.980 29.850 885.360 30.230 ;
        RECT 890.690 30.150 892.430 30.440 ;
        RECT 894.480 30.100 895.680 30.390 ;
        RECT 897.190 30.060 899.820 30.515 ;
        RECT 901.400 30.165 901.780 30.545 ;
        RECT 806.135 29.400 819.960 29.700 ;
        RECT 821.635 29.235 837.645 29.610 ;
        RECT 855.570 29.225 876.345 29.600 ;
        RECT 806.140 28.655 824.560 28.955 ;
        RECT 826.005 28.645 853.315 28.985 ;
        RECT 805.620 27.940 812.880 28.240 ;
        RECT 625.295 27.515 643.965 27.525 ;
        RECT 625.295 27.505 682.665 27.515 ;
        RECT 625.295 27.205 691.670 27.505 ;
        RECT 790.675 27.320 794.800 27.590 ;
        RECT 806.175 27.405 810.260 27.675 ;
        RECT 816.580 27.640 820.330 27.915 ;
        RECT 821.635 27.880 847.865 28.270 ;
        RECT 854.600 27.870 886.565 28.260 ;
        RECT 899.375 27.630 902.505 27.905 ;
        RECT 903.250 27.870 903.630 35.030 ;
        RECT 952.880 32.925 954.080 33.305 ;
        RECT 904.490 32.570 911.230 32.870 ;
        RECT 955.835 32.710 958.110 33.220 ;
        RECT 960.735 32.710 963.035 33.220 ;
        RECT 965.330 32.710 967.610 33.220 ;
        RECT 972.405 33.025 973.640 33.405 ;
        RECT 905.080 30.775 908.535 31.215 ;
        RECT 908.825 30.575 909.205 30.955 ;
        RECT 911.540 30.615 911.920 30.995 ;
        RECT 915.725 30.565 916.105 30.945 ;
        RECT 952.880 30.625 956.140 31.005 ;
        RECT 956.880 30.625 960.140 31.005 ;
        RECT 966.380 30.625 969.640 31.005 ;
        RECT 970.380 30.625 973.640 31.005 ;
        RECT 906.150 30.150 907.890 30.440 ;
        RECT 909.940 30.100 911.140 30.390 ;
        RECT 912.650 30.070 915.275 30.480 ;
        RECT 916.860 30.165 917.240 30.545 ;
        RECT 903.895 29.390 919.815 29.690 ;
        RECT 953.545 28.975 975.830 29.050 ;
        RECT 904.430 28.645 921.375 28.945 ;
        RECT 953.545 28.710 979.890 28.975 ;
        RECT 975.715 28.635 979.890 28.710 ;
        RECT 914.835 27.630 922.535 27.905 ;
        RECT 985.875 27.880 986.255 35.040 ;
        RECT 987.705 30.825 991.080 31.225 ;
        RECT 991.450 30.585 991.830 30.965 ;
        RECT 994.165 30.625 994.545 31.005 ;
        RECT 998.350 30.575 998.730 30.955 ;
        RECT 988.775 30.160 990.515 30.450 ;
        RECT 992.565 30.110 993.765 30.400 ;
        RECT 995.275 30.080 997.885 30.505 ;
        RECT 999.485 30.175 999.865 30.555 ;
        RECT 987.020 29.400 1000.585 29.715 ;
        RECT 987.015 28.655 1000.575 28.955 ;
        RECT 987.035 27.940 993.760 28.240 ;
        RECT 997.460 27.640 1000.565 27.915 ;
        RECT 1001.335 27.880 1001.715 35.040 ;
        RECT 1057.895 35.030 1114.250 35.040 ;
        RECT 1017.975 34.045 1055.525 34.055 ;
        RECT 1017.975 33.770 1083.655 34.045 ;
        RECT 1054.880 33.760 1083.655 33.770 ;
        RECT 1085.325 33.740 1092.030 34.040 ;
        RECT 1019.485 32.860 1020.940 33.240 ;
        RECT 1021.680 32.860 1022.880 33.240 ;
        RECT 1024.635 32.645 1026.910 33.155 ;
        RECT 1029.535 32.645 1031.835 33.155 ;
        RECT 1034.130 32.645 1036.410 33.155 ;
        RECT 1041.205 32.960 1042.440 33.340 ;
        RECT 1043.180 32.960 1044.460 33.340 ;
        RECT 1058.185 32.850 1059.640 33.230 ;
        RECT 1042.620 32.605 1043.000 32.640 ;
        RECT 1063.335 32.635 1065.610 33.145 ;
        RECT 1068.235 32.635 1070.535 33.145 ;
        RECT 1072.830 32.635 1075.110 33.145 ;
        RECT 1081.880 32.950 1083.160 33.330 ;
        RECT 1021.120 32.500 1021.500 32.540 ;
        RECT 1021.050 32.195 1023.885 32.500 ;
        RECT 1039.865 32.295 1043.000 32.605 ;
        RECT 1081.320 32.595 1081.700 32.630 ;
        RECT 1059.820 32.490 1060.200 32.530 ;
        RECT 1042.620 32.260 1043.000 32.295 ;
        RECT 1021.120 32.160 1021.500 32.195 ;
        RECT 1059.750 32.185 1062.585 32.490 ;
        RECT 1078.565 32.285 1081.700 32.595 ;
        RECT 1081.320 32.250 1081.700 32.285 ;
        RECT 1059.820 32.150 1060.200 32.185 ;
        RECT 1003.165 30.785 1006.570 31.225 ;
        RECT 1006.910 30.585 1007.290 30.965 ;
        RECT 1009.625 30.625 1010.005 31.005 ;
        RECT 1013.810 30.575 1014.190 30.955 ;
        RECT 1019.645 30.560 1020.940 30.940 ;
        RECT 1021.680 30.560 1024.940 30.940 ;
        RECT 1025.680 30.560 1028.940 30.940 ;
        RECT 1029.680 30.560 1030.865 30.940 ;
        RECT 1033.130 30.560 1034.440 30.940 ;
        RECT 1035.180 30.560 1038.440 30.940 ;
        RECT 1039.180 30.560 1042.440 30.940 ;
        RECT 1043.180 30.560 1044.195 30.940 ;
        RECT 1004.235 30.160 1005.975 30.450 ;
        RECT 1008.025 30.110 1009.225 30.400 ;
        RECT 1010.735 30.080 1013.330 30.455 ;
        RECT 1014.945 30.175 1015.325 30.555 ;
        RECT 1058.345 30.550 1059.640 30.930 ;
        RECT 1064.380 30.550 1067.640 30.930 ;
        RECT 1068.380 30.550 1069.565 30.930 ;
        RECT 1071.830 30.550 1073.140 30.930 ;
        RECT 1073.880 30.550 1077.140 30.930 ;
        RECT 1081.880 30.550 1082.895 30.930 ;
        RECT 1085.960 30.795 1089.375 31.215 ;
        RECT 1089.705 30.575 1090.085 30.955 ;
        RECT 1092.420 30.615 1092.800 30.995 ;
        RECT 1096.605 30.565 1096.985 30.945 ;
        RECT 1021.120 29.860 1021.500 30.240 ;
        RECT 1025.120 29.860 1025.500 30.240 ;
        RECT 1029.120 30.195 1029.500 30.240 ;
        RECT 1034.620 30.195 1035.000 30.240 ;
        RECT 1029.070 29.880 1035.005 30.195 ;
        RECT 1029.120 29.860 1029.500 29.880 ;
        RECT 1034.620 29.860 1035.000 29.880 ;
        RECT 1038.620 29.860 1039.000 30.240 ;
        RECT 1042.620 29.860 1043.000 30.240 ;
        RECT 1059.820 29.850 1060.200 30.230 ;
        RECT 1063.820 29.850 1064.200 30.230 ;
        RECT 1067.820 30.185 1068.200 30.230 ;
        RECT 1073.320 30.185 1073.700 30.230 ;
        RECT 1067.770 29.870 1073.705 30.185 ;
        RECT 1067.820 29.850 1068.200 29.870 ;
        RECT 1073.320 29.850 1073.700 29.870 ;
        RECT 1077.320 29.850 1077.700 30.230 ;
        RECT 1081.320 29.850 1081.700 30.230 ;
        RECT 1087.030 30.150 1088.770 30.440 ;
        RECT 1090.820 30.100 1092.020 30.390 ;
        RECT 1093.530 30.060 1096.160 30.515 ;
        RECT 1097.740 30.165 1098.120 30.545 ;
        RECT 1002.475 29.400 1016.300 29.700 ;
        RECT 1017.975 29.235 1033.985 29.610 ;
        RECT 1051.910 29.225 1072.685 29.600 ;
        RECT 1002.480 28.655 1020.900 28.955 ;
        RECT 1022.345 28.645 1049.655 28.985 ;
        RECT 1001.960 27.940 1009.220 28.240 ;
        RECT 821.635 27.515 840.305 27.525 ;
        RECT 821.635 27.505 879.005 27.515 ;
        RECT 821.635 27.205 888.010 27.505 ;
        RECT 987.015 27.320 991.140 27.590 ;
        RECT 1002.515 27.405 1006.600 27.675 ;
        RECT 1012.920 27.640 1016.670 27.915 ;
        RECT 1017.975 27.880 1044.205 28.270 ;
        RECT 1050.940 27.870 1082.905 28.260 ;
        RECT 1095.715 27.630 1098.845 27.905 ;
        RECT 1099.590 27.870 1099.970 35.030 ;
        RECT 1149.205 32.930 1150.405 33.310 ;
        RECT 1100.830 32.570 1107.570 32.870 ;
        RECT 1152.160 32.715 1154.435 33.225 ;
        RECT 1157.060 32.715 1159.360 33.225 ;
        RECT 1161.655 32.715 1163.935 33.225 ;
        RECT 1168.730 33.030 1169.965 33.410 ;
        RECT 1101.420 30.775 1104.875 31.215 ;
        RECT 1105.165 30.575 1105.545 30.955 ;
        RECT 1107.880 30.615 1108.260 30.995 ;
        RECT 1112.065 30.565 1112.445 30.945 ;
        RECT 1149.205 30.630 1152.465 31.010 ;
        RECT 1153.205 30.630 1156.465 31.010 ;
        RECT 1162.705 30.630 1165.965 31.010 ;
        RECT 1166.705 30.630 1169.965 31.010 ;
        RECT 1102.490 30.150 1104.230 30.440 ;
        RECT 1106.280 30.100 1107.480 30.390 ;
        RECT 1108.990 30.070 1111.615 30.480 ;
        RECT 1113.200 30.165 1113.580 30.545 ;
        RECT 1100.235 29.390 1116.155 29.690 ;
        RECT 1149.870 28.980 1172.155 29.055 ;
        RECT 1100.770 28.645 1117.715 28.945 ;
        RECT 1149.870 28.715 1176.215 28.980 ;
        RECT 1172.040 28.640 1176.215 28.715 ;
        RECT 1111.175 27.630 1118.875 27.905 ;
        RECT 1182.215 27.880 1182.595 35.040 ;
        RECT 1184.045 30.825 1187.420 31.225 ;
        RECT 1187.790 30.585 1188.170 30.965 ;
        RECT 1190.505 30.625 1190.885 31.005 ;
        RECT 1194.690 30.575 1195.070 30.955 ;
        RECT 1185.115 30.160 1186.855 30.450 ;
        RECT 1188.905 30.110 1190.105 30.400 ;
        RECT 1191.615 30.080 1194.225 30.505 ;
        RECT 1195.825 30.175 1196.205 30.555 ;
        RECT 1183.360 29.400 1196.925 29.715 ;
        RECT 1183.355 28.655 1196.915 28.955 ;
        RECT 1183.375 27.940 1190.100 28.240 ;
        RECT 1193.800 27.640 1196.905 27.915 ;
        RECT 1197.675 27.880 1198.055 35.040 ;
        RECT 1254.235 35.030 1310.590 35.040 ;
        RECT 1214.315 34.045 1251.865 34.055 ;
        RECT 1214.315 33.770 1279.995 34.045 ;
        RECT 1251.220 33.760 1279.995 33.770 ;
        RECT 1281.665 33.740 1288.370 34.040 ;
        RECT 1215.825 32.860 1217.280 33.240 ;
        RECT 1218.020 32.860 1219.220 33.240 ;
        RECT 1220.975 32.645 1223.250 33.155 ;
        RECT 1225.875 32.645 1228.175 33.155 ;
        RECT 1230.470 32.645 1232.750 33.155 ;
        RECT 1237.545 32.960 1238.780 33.340 ;
        RECT 1239.520 32.960 1240.800 33.340 ;
        RECT 1254.525 32.850 1255.980 33.230 ;
        RECT 1256.720 32.850 1257.920 33.230 ;
        RECT 1238.960 32.605 1239.340 32.640 ;
        RECT 1259.675 32.635 1261.950 33.145 ;
        RECT 1264.575 32.635 1266.875 33.145 ;
        RECT 1269.170 32.635 1271.450 33.145 ;
        RECT 1276.245 32.950 1277.480 33.330 ;
        RECT 1278.220 32.950 1279.500 33.330 ;
        RECT 1217.460 32.500 1217.840 32.540 ;
        RECT 1217.390 32.195 1220.225 32.500 ;
        RECT 1236.205 32.295 1239.340 32.605 ;
        RECT 1277.660 32.595 1278.040 32.630 ;
        RECT 1256.160 32.490 1256.540 32.530 ;
        RECT 1238.960 32.260 1239.340 32.295 ;
        RECT 1217.460 32.160 1217.840 32.195 ;
        RECT 1256.090 32.185 1258.925 32.490 ;
        RECT 1274.905 32.285 1278.040 32.595 ;
        RECT 1277.660 32.250 1278.040 32.285 ;
        RECT 1256.160 32.150 1256.540 32.185 ;
        RECT 1199.505 30.785 1202.910 31.225 ;
        RECT 1203.250 30.585 1203.630 30.965 ;
        RECT 1205.965 30.625 1206.345 31.005 ;
        RECT 1210.150 30.575 1210.530 30.955 ;
        RECT 1215.985 30.560 1217.280 30.940 ;
        RECT 1218.020 30.560 1221.280 30.940 ;
        RECT 1222.020 30.560 1225.280 30.940 ;
        RECT 1226.020 30.560 1227.205 30.940 ;
        RECT 1229.470 30.560 1230.780 30.940 ;
        RECT 1231.520 30.560 1234.780 30.940 ;
        RECT 1235.520 30.560 1238.780 30.940 ;
        RECT 1239.520 30.560 1240.535 30.940 ;
        RECT 1200.575 30.160 1202.315 30.450 ;
        RECT 1204.365 30.110 1205.565 30.400 ;
        RECT 1207.075 30.080 1209.670 30.455 ;
        RECT 1211.285 30.175 1211.665 30.555 ;
        RECT 1254.685 30.550 1255.980 30.930 ;
        RECT 1256.720 30.550 1259.980 30.930 ;
        RECT 1260.720 30.550 1263.980 30.930 ;
        RECT 1264.720 30.550 1265.905 30.930 ;
        RECT 1268.170 30.550 1269.480 30.930 ;
        RECT 1270.220 30.550 1273.480 30.930 ;
        RECT 1274.220 30.550 1277.480 30.930 ;
        RECT 1278.220 30.550 1279.235 30.930 ;
        RECT 1282.300 30.795 1285.715 31.215 ;
        RECT 1286.045 30.575 1286.425 30.955 ;
        RECT 1288.760 30.615 1289.140 30.995 ;
        RECT 1292.945 30.565 1293.325 30.945 ;
        RECT 1217.460 29.860 1217.840 30.240 ;
        RECT 1221.460 29.860 1221.840 30.240 ;
        RECT 1225.460 30.195 1225.840 30.240 ;
        RECT 1230.960 30.195 1231.340 30.240 ;
        RECT 1225.410 29.880 1231.345 30.195 ;
        RECT 1225.460 29.860 1225.840 29.880 ;
        RECT 1230.960 29.860 1231.340 29.880 ;
        RECT 1234.960 29.860 1235.340 30.240 ;
        RECT 1238.960 29.860 1239.340 30.240 ;
        RECT 1256.160 29.850 1256.540 30.230 ;
        RECT 1260.160 29.850 1260.540 30.230 ;
        RECT 1264.160 30.185 1264.540 30.230 ;
        RECT 1269.660 30.185 1270.040 30.230 ;
        RECT 1264.110 29.870 1270.045 30.185 ;
        RECT 1264.160 29.850 1264.540 29.870 ;
        RECT 1269.660 29.850 1270.040 29.870 ;
        RECT 1273.660 29.850 1274.040 30.230 ;
        RECT 1277.660 29.850 1278.040 30.230 ;
        RECT 1283.370 30.150 1285.110 30.440 ;
        RECT 1287.160 30.100 1288.360 30.390 ;
        RECT 1289.870 30.060 1292.500 30.515 ;
        RECT 1294.080 30.165 1294.460 30.545 ;
        RECT 1198.815 29.400 1212.640 29.700 ;
        RECT 1214.315 29.235 1230.325 29.610 ;
        RECT 1248.250 29.225 1269.025 29.600 ;
        RECT 1281.650 29.390 1295.265 29.690 ;
        RECT 1198.820 28.655 1217.240 28.955 ;
        RECT 1218.685 28.645 1245.995 28.985 ;
        RECT 1257.385 28.635 1279.940 28.975 ;
        RECT 1281.050 28.645 1295.695 28.945 ;
        RECT 1198.300 27.940 1205.560 28.240 ;
        RECT 1017.975 27.515 1036.645 27.525 ;
        RECT 1017.975 27.505 1075.345 27.515 ;
        RECT 1017.975 27.205 1084.350 27.505 ;
        RECT 1183.355 27.320 1187.480 27.590 ;
        RECT 1198.855 27.405 1202.940 27.675 ;
        RECT 1209.260 27.640 1213.010 27.915 ;
        RECT 1214.315 27.880 1240.545 28.270 ;
        RECT 1247.280 27.870 1279.245 28.260 ;
        RECT 1292.055 27.630 1295.185 27.905 ;
        RECT 1295.930 27.870 1296.310 35.030 ;
        RECT 1297.170 32.570 1303.910 32.870 ;
        RECT 1297.760 30.775 1301.215 31.215 ;
        RECT 1304.220 30.615 1304.600 30.995 ;
        RECT 1302.620 30.100 1303.820 30.390 ;
        RECT 1309.540 30.165 1309.920 30.545 ;
        RECT 1296.575 29.390 1312.495 29.690 ;
        RECT 1297.110 28.645 1314.055 28.945 ;
        RECT 1214.315 27.515 1232.985 27.525 ;
        RECT 1214.315 27.505 1271.685 27.515 ;
        RECT 1214.315 27.205 1280.690 27.505 ;
        RECT 655.105 27.195 691.670 27.205 ;
        RECT 851.445 27.195 888.010 27.205 ;
        RECT 1047.785 27.195 1084.350 27.205 ;
        RECT 1244.125 27.195 1280.690 27.205 ;
        RECT 458.730 27.160 495.295 27.170 ;
        RECT -59.660 25.925 -56.095 25.935 ;
        RECT -59.660 25.600 -55.300 25.925 ;
        RECT -56.255 25.590 -55.300 25.600 ;
        RECT -79.065 24.960 -75.765 25.340 ;
        RECT -75.065 24.960 -71.765 25.340 ;
        RECT -65.565 24.960 -62.265 25.340 ;
        RECT -61.565 24.960 -58.265 25.340 ;
        RECT -79.065 22.960 -77.780 23.340 ;
        RECT -59.750 22.960 -58.265 23.340 ;
        RECT -77.560 22.280 -76.040 22.640 ;
        RECT 4.055 20.930 4.435 26.760 ;
        RECT 8.895 26.160 15.285 26.450 ;
        RECT 8.310 25.580 18.965 25.915 ;
        RECT 5.875 24.245 6.255 24.625 ;
        RECT 8.280 24.260 10.060 24.550 ;
        RECT 11.535 24.350 12.725 24.635 ;
        RECT 15.655 24.230 16.965 24.550 ;
        RECT 7.010 23.645 7.390 24.025 ;
        RECT 10.755 23.685 11.135 24.065 ;
        RECT 13.465 23.675 13.845 24.055 ;
        RECT 14.875 23.520 18.055 23.840 ;
        RECT 4.805 20.930 8.900 20.935 ;
        RECT 19.515 20.930 19.895 26.760 ;
        RECT 120.145 26.750 124.275 27.050 ;
        RECT 35.625 26.540 71.535 26.550 ;
        RECT 24.355 26.160 30.745 26.450 ;
        RECT 35.625 26.280 102.930 26.540 ;
        RECT 71.185 26.270 102.930 26.280 ;
        RECT 107.150 26.150 113.540 26.440 ;
        RECT 23.770 25.580 34.275 25.915 ;
        RECT 59.245 25.715 69.795 26.050 ;
        RECT 106.565 25.570 117.045 25.905 ;
        RECT 39.840 25.075 43.140 25.455 ;
        RECT 43.840 25.075 47.140 25.455 ;
        RECT 53.340 25.075 56.640 25.455 ;
        RECT 57.340 25.075 60.640 25.455 ;
        RECT 76.535 25.065 77.840 25.445 ;
        RECT 82.540 25.065 85.840 25.445 ;
        RECT 86.540 25.065 87.900 25.445 ;
        RECT 89.875 25.065 91.340 25.445 ;
        RECT 92.040 25.065 95.340 25.445 ;
        RECT 100.040 25.065 101.220 25.445 ;
        RECT 39.300 24.730 39.680 24.765 ;
        RECT 21.335 24.245 21.715 24.625 ;
        RECT 23.740 24.260 25.520 24.550 ;
        RECT 26.995 24.350 28.185 24.635 ;
        RECT 31.115 24.230 32.425 24.550 ;
        RECT 39.035 24.420 42.045 24.730 ;
        RECT 39.300 24.385 39.680 24.420 ;
        RECT 43.300 24.385 44.390 24.765 ;
        RECT 47.300 24.760 47.680 24.765 ;
        RECT 44.820 24.395 47.685 24.760 ;
        RECT 52.800 24.740 53.180 24.765 ;
        RECT 52.785 24.420 54.930 24.740 ;
        RECT 47.300 24.385 47.680 24.395 ;
        RECT 52.800 24.385 53.180 24.420 ;
        RECT 55.845 24.385 57.180 24.765 ;
        RECT 60.800 24.745 61.180 24.765 ;
        RECT 58.335 24.425 61.245 24.745 ;
        RECT 78.000 24.720 78.380 24.755 ;
        RECT 60.800 24.385 61.180 24.425 ;
        RECT 77.735 24.410 80.745 24.720 ;
        RECT 78.000 24.375 78.380 24.410 ;
        RECT 82.000 24.375 83.090 24.755 ;
        RECT 86.000 24.750 86.380 24.755 ;
        RECT 83.520 24.385 86.385 24.750 ;
        RECT 91.500 24.730 91.880 24.755 ;
        RECT 91.485 24.410 93.630 24.730 ;
        RECT 86.000 24.375 86.380 24.385 ;
        RECT 91.500 24.375 91.880 24.410 ;
        RECT 94.545 24.375 95.880 24.755 ;
        RECT 99.500 24.735 99.880 24.755 ;
        RECT 97.035 24.415 99.945 24.735 ;
        RECT 99.500 24.375 99.880 24.415 ;
        RECT 104.130 24.235 104.510 24.615 ;
        RECT 106.535 24.250 108.315 24.540 ;
        RECT 109.790 24.340 110.980 24.625 ;
        RECT 113.910 24.220 115.220 24.540 ;
        RECT 22.470 23.645 22.850 24.025 ;
        RECT 26.215 23.685 26.595 24.065 ;
        RECT 28.925 23.675 29.305 24.055 ;
        RECT 30.335 23.520 33.515 23.840 ;
        RECT 105.265 23.635 105.645 24.015 ;
        RECT 109.010 23.675 109.390 24.055 ;
        RECT 111.720 23.665 112.100 24.045 ;
        RECT 113.130 23.510 116.310 23.830 ;
        RECT 39.840 23.075 41.125 23.455 ;
        RECT 59.155 23.075 60.640 23.455 ;
        RECT 76.350 23.065 77.840 23.445 ;
        RECT 100.040 23.065 101.115 23.445 ;
        RECT 39.300 22.385 40.390 22.765 ;
        RECT 41.345 22.395 42.865 22.755 ;
        RECT 43.785 22.390 56.635 22.725 ;
        RECT 60.800 22.720 61.180 22.765 ;
        RECT 60.065 22.420 61.375 22.720 ;
        RECT 60.800 22.385 61.180 22.420 ;
        RECT 78.000 22.375 79.090 22.755 ;
        RECT 80.045 22.385 81.565 22.745 ;
        RECT 82.485 22.380 95.335 22.715 ;
        RECT 99.500 22.710 99.880 22.755 ;
        RECT 98.765 22.410 100.075 22.710 ;
        RECT 99.500 22.375 99.880 22.410 ;
        RECT 68.560 21.875 101.510 21.880 ;
        RECT 36.155 21.525 101.510 21.875 ;
        RECT 68.560 21.515 101.510 21.525 ;
        RECT 103.305 21.505 107.565 21.860 ;
        RECT 20.265 20.930 24.360 20.935 ;
        RECT 3.685 20.925 8.900 20.930 ;
        RECT 19.145 20.925 24.360 20.930 ;
        RECT 34.605 20.925 74.855 20.930 ;
        RECT 3.685 20.920 74.855 20.925 ;
        RECT 101.510 20.920 107.155 20.925 ;
        RECT 117.770 20.920 118.150 26.750 ;
        RECT 126.650 26.700 131.150 27.010 ;
        RECT 202.795 26.760 206.925 27.060 ;
        RECT 122.610 26.150 129.000 26.440 ;
        RECT 122.025 25.570 138.045 25.905 ;
        RECT 186.805 25.770 192.775 26.105 ;
        RECT 121.375 24.985 124.295 25.285 ;
        RECT 127.840 24.970 131.210 25.270 ;
        RECT 167.400 25.130 170.700 25.510 ;
        RECT 171.400 25.130 174.700 25.510 ;
        RECT 180.900 25.130 184.200 25.510 ;
        RECT 184.900 25.130 188.200 25.510 ;
        RECT 119.590 24.235 119.970 24.615 ;
        RECT 121.995 24.250 123.775 24.540 ;
        RECT 125.250 24.340 126.440 24.625 ;
        RECT 129.370 24.220 130.680 24.540 ;
        RECT 120.725 23.635 121.105 24.015 ;
        RECT 124.470 23.675 124.850 24.055 ;
        RECT 127.180 23.665 127.560 24.045 ;
        RECT 128.590 23.510 131.770 23.830 ;
        RECT 167.400 23.130 168.685 23.510 ;
        RECT 186.715 23.130 188.200 23.510 ;
        RECT 118.870 22.425 123.020 22.695 ;
        RECT 168.905 22.450 170.425 22.810 ;
        RECT 118.520 20.920 122.615 20.925 ;
        RECT 3.685 20.915 107.155 20.920 ;
        RECT 117.400 20.915 122.615 20.920 ;
        RECT -82.750 19.915 -56.095 20.815 ;
        RECT 3.685 20.030 132.430 20.915 ;
        RECT 163.715 20.085 190.370 20.985 ;
        RECT 200.420 20.930 200.800 26.760 ;
        RECT 209.300 26.710 213.800 27.020 ;
        RECT 218.255 26.760 222.385 27.060 ;
        RECT 205.260 26.160 211.650 26.450 ;
        RECT 204.675 25.580 215.330 25.915 ;
        RECT 204.025 24.995 206.945 25.295 ;
        RECT 210.490 24.980 213.860 25.280 ;
        RECT 202.240 24.245 202.620 24.625 ;
        RECT 204.645 24.260 206.425 24.550 ;
        RECT 207.900 24.350 209.090 24.635 ;
        RECT 212.020 24.230 213.330 24.550 ;
        RECT 203.375 23.645 203.755 24.025 ;
        RECT 207.120 23.685 207.500 24.065 ;
        RECT 209.830 23.675 210.210 24.055 ;
        RECT 211.240 23.520 214.420 23.840 ;
        RECT 201.170 20.930 205.265 20.935 ;
        RECT 215.880 20.930 216.260 26.760 ;
        RECT 224.760 26.710 229.260 27.020 ;
        RECT 316.510 26.750 320.640 27.050 ;
        RECT 231.990 26.540 267.900 26.550 ;
        RECT 220.720 26.160 227.110 26.450 ;
        RECT 231.990 26.280 299.295 26.540 ;
        RECT 267.550 26.270 299.295 26.280 ;
        RECT 303.515 26.150 309.905 26.440 ;
        RECT 220.135 25.580 230.640 25.915 ;
        RECT 255.610 25.715 266.160 26.050 ;
        RECT 302.930 25.570 313.410 25.905 ;
        RECT 219.485 24.995 222.405 25.295 ;
        RECT 225.950 24.980 229.320 25.280 ;
        RECT 234.200 25.075 235.505 25.455 ;
        RECT 236.205 25.075 239.505 25.455 ;
        RECT 240.205 25.075 243.505 25.455 ;
        RECT 244.205 25.075 245.565 25.455 ;
        RECT 247.540 25.075 249.005 25.455 ;
        RECT 249.705 25.075 253.005 25.455 ;
        RECT 253.705 25.075 257.005 25.455 ;
        RECT 257.705 25.075 258.885 25.455 ;
        RECT 272.900 25.065 274.205 25.445 ;
        RECT 278.905 25.065 282.205 25.445 ;
        RECT 282.905 25.065 284.265 25.445 ;
        RECT 286.240 25.065 287.705 25.445 ;
        RECT 288.405 25.065 291.705 25.445 ;
        RECT 296.405 25.065 297.585 25.445 ;
        RECT 235.665 24.730 236.045 24.765 ;
        RECT 217.700 24.245 218.080 24.625 ;
        RECT 220.105 24.260 221.885 24.550 ;
        RECT 223.360 24.350 224.550 24.635 ;
        RECT 227.480 24.230 228.790 24.550 ;
        RECT 235.400 24.420 238.410 24.730 ;
        RECT 235.665 24.385 236.045 24.420 ;
        RECT 239.665 24.385 240.755 24.765 ;
        RECT 243.665 24.760 244.045 24.765 ;
        RECT 241.185 24.395 244.050 24.760 ;
        RECT 249.165 24.740 249.545 24.765 ;
        RECT 249.150 24.420 251.295 24.740 ;
        RECT 243.665 24.385 244.045 24.395 ;
        RECT 249.165 24.385 249.545 24.420 ;
        RECT 252.210 24.385 253.545 24.765 ;
        RECT 257.165 24.745 257.545 24.765 ;
        RECT 254.700 24.425 257.610 24.745 ;
        RECT 274.365 24.720 274.745 24.755 ;
        RECT 257.165 24.385 257.545 24.425 ;
        RECT 274.100 24.410 277.110 24.720 ;
        RECT 274.365 24.375 274.745 24.410 ;
        RECT 278.365 24.375 279.455 24.755 ;
        RECT 282.365 24.750 282.745 24.755 ;
        RECT 279.885 24.385 282.750 24.750 ;
        RECT 287.865 24.730 288.245 24.755 ;
        RECT 287.850 24.410 289.995 24.730 ;
        RECT 282.365 24.375 282.745 24.385 ;
        RECT 287.865 24.375 288.245 24.410 ;
        RECT 290.910 24.375 292.245 24.755 ;
        RECT 295.865 24.735 296.245 24.755 ;
        RECT 293.400 24.415 296.310 24.735 ;
        RECT 295.865 24.375 296.245 24.415 ;
        RECT 300.495 24.235 300.875 24.615 ;
        RECT 302.900 24.250 304.680 24.540 ;
        RECT 306.155 24.340 307.345 24.625 ;
        RECT 310.275 24.220 311.585 24.540 ;
        RECT 218.835 23.645 219.215 24.025 ;
        RECT 222.580 23.685 222.960 24.065 ;
        RECT 225.290 23.675 225.670 24.055 ;
        RECT 226.700 23.520 229.880 23.840 ;
        RECT 301.630 23.635 302.010 24.015 ;
        RECT 305.375 23.675 305.755 24.055 ;
        RECT 308.085 23.665 308.465 24.045 ;
        RECT 309.495 23.510 312.675 23.830 ;
        RECT 234.015 23.075 235.505 23.455 ;
        RECT 236.205 23.075 237.490 23.455 ;
        RECT 255.520 23.075 257.005 23.455 ;
        RECT 257.705 23.075 258.780 23.455 ;
        RECT 272.715 23.065 274.205 23.445 ;
        RECT 296.405 23.065 297.480 23.445 ;
        RECT 235.665 22.385 236.755 22.765 ;
        RECT 237.710 22.395 239.230 22.755 ;
        RECT 240.150 22.390 253.000 22.725 ;
        RECT 257.165 22.720 257.545 22.765 ;
        RECT 256.430 22.420 257.740 22.720 ;
        RECT 257.165 22.385 257.545 22.420 ;
        RECT 274.365 22.375 275.455 22.755 ;
        RECT 276.410 22.385 277.930 22.745 ;
        RECT 278.850 22.380 291.700 22.715 ;
        RECT 295.865 22.710 296.245 22.755 ;
        RECT 295.130 22.410 296.440 22.710 ;
        RECT 295.865 22.375 296.245 22.410 ;
        RECT 264.925 21.875 297.875 21.880 ;
        RECT 232.520 21.525 297.875 21.875 ;
        RECT 264.925 21.515 297.875 21.525 ;
        RECT 299.670 21.505 303.930 21.860 ;
        RECT 216.630 20.930 220.725 20.935 ;
        RECT 200.050 20.925 205.265 20.930 ;
        RECT 215.510 20.925 220.725 20.930 ;
        RECT 230.970 20.925 271.220 20.930 ;
        RECT 200.050 20.920 271.220 20.925 ;
        RECT 297.875 20.920 303.520 20.925 ;
        RECT 314.135 20.920 314.515 26.750 ;
        RECT 323.015 26.700 327.515 27.010 ;
        RECT 399.195 26.710 403.325 27.010 ;
        RECT 318.975 26.150 325.365 26.440 ;
        RECT 318.390 25.570 334.410 25.905 ;
        RECT 383.195 25.730 389.165 26.065 ;
        RECT 317.740 24.985 320.660 25.285 ;
        RECT 324.205 24.970 327.575 25.270 ;
        RECT 363.790 25.090 367.090 25.470 ;
        RECT 367.790 25.090 371.090 25.470 ;
        RECT 377.290 25.090 380.590 25.470 ;
        RECT 381.290 25.090 384.590 25.470 ;
        RECT 315.955 24.235 316.335 24.615 ;
        RECT 318.360 24.250 320.140 24.540 ;
        RECT 321.615 24.340 322.805 24.625 ;
        RECT 325.735 24.220 327.045 24.540 ;
        RECT 317.090 23.635 317.470 24.015 ;
        RECT 320.835 23.675 321.215 24.055 ;
        RECT 323.545 23.665 323.925 24.045 ;
        RECT 324.955 23.510 328.135 23.830 ;
        RECT 363.790 23.090 365.075 23.470 ;
        RECT 383.105 23.090 384.590 23.470 ;
        RECT 315.235 22.425 319.385 22.695 ;
        RECT 365.295 22.410 366.815 22.770 ;
        RECT 314.885 20.920 318.980 20.925 ;
        RECT 200.050 20.915 303.520 20.920 ;
        RECT 313.765 20.915 318.980 20.920 ;
        RECT 200.050 20.030 328.795 20.915 ;
        RECT 360.105 20.045 386.760 20.945 ;
        RECT 396.820 20.880 397.200 26.710 ;
        RECT 405.700 26.660 410.200 26.970 ;
        RECT 414.655 26.710 418.785 27.010 ;
        RECT 401.660 26.110 408.050 26.400 ;
        RECT 401.075 25.530 411.730 25.865 ;
        RECT 400.425 24.945 403.345 25.245 ;
        RECT 406.890 24.930 410.260 25.230 ;
        RECT 398.640 24.195 399.020 24.575 ;
        RECT 401.045 24.210 402.825 24.500 ;
        RECT 404.300 24.300 405.490 24.585 ;
        RECT 408.420 24.180 409.730 24.500 ;
        RECT 399.775 23.595 400.155 23.975 ;
        RECT 403.520 23.635 403.900 24.015 ;
        RECT 406.230 23.625 406.610 24.005 ;
        RECT 407.640 23.470 410.820 23.790 ;
        RECT 397.570 20.880 401.665 20.885 ;
        RECT 412.280 20.880 412.660 26.710 ;
        RECT 421.160 26.660 425.660 26.970 ;
        RECT 512.910 26.700 517.040 27.000 ;
        RECT 428.390 26.490 464.300 26.500 ;
        RECT 417.120 26.110 423.510 26.400 ;
        RECT 428.390 26.230 495.695 26.490 ;
        RECT 463.950 26.220 495.695 26.230 ;
        RECT 499.915 26.100 506.305 26.390 ;
        RECT 416.535 25.530 427.040 25.865 ;
        RECT 452.010 25.665 462.560 26.000 ;
        RECT 499.330 25.520 509.810 25.855 ;
        RECT 415.885 24.945 418.805 25.245 ;
        RECT 422.350 24.930 425.720 25.230 ;
        RECT 430.600 25.025 431.905 25.405 ;
        RECT 432.605 25.025 435.905 25.405 ;
        RECT 436.605 25.025 439.905 25.405 ;
        RECT 440.605 25.025 441.965 25.405 ;
        RECT 443.940 25.025 445.405 25.405 ;
        RECT 446.105 25.025 449.405 25.405 ;
        RECT 450.105 25.025 453.405 25.405 ;
        RECT 454.105 25.025 455.285 25.405 ;
        RECT 469.300 25.015 470.605 25.395 ;
        RECT 475.305 25.015 478.605 25.395 ;
        RECT 479.305 25.015 480.665 25.395 ;
        RECT 482.640 25.015 484.105 25.395 ;
        RECT 484.805 25.015 488.105 25.395 ;
        RECT 492.805 25.015 493.985 25.395 ;
        RECT 432.065 24.680 432.445 24.715 ;
        RECT 414.100 24.195 414.480 24.575 ;
        RECT 416.505 24.210 418.285 24.500 ;
        RECT 419.760 24.300 420.950 24.585 ;
        RECT 423.880 24.180 425.190 24.500 ;
        RECT 431.800 24.370 434.810 24.680 ;
        RECT 432.065 24.335 432.445 24.370 ;
        RECT 436.065 24.335 437.155 24.715 ;
        RECT 440.065 24.710 440.445 24.715 ;
        RECT 437.585 24.345 440.450 24.710 ;
        RECT 445.565 24.690 445.945 24.715 ;
        RECT 445.550 24.370 447.695 24.690 ;
        RECT 440.065 24.335 440.445 24.345 ;
        RECT 445.565 24.335 445.945 24.370 ;
        RECT 448.610 24.335 449.945 24.715 ;
        RECT 453.565 24.695 453.945 24.715 ;
        RECT 451.100 24.375 454.010 24.695 ;
        RECT 470.765 24.670 471.145 24.705 ;
        RECT 453.565 24.335 453.945 24.375 ;
        RECT 470.500 24.360 473.510 24.670 ;
        RECT 470.765 24.325 471.145 24.360 ;
        RECT 474.765 24.325 475.855 24.705 ;
        RECT 478.765 24.700 479.145 24.705 ;
        RECT 476.285 24.335 479.150 24.700 ;
        RECT 484.265 24.680 484.645 24.705 ;
        RECT 484.250 24.360 486.395 24.680 ;
        RECT 478.765 24.325 479.145 24.335 ;
        RECT 484.265 24.325 484.645 24.360 ;
        RECT 487.310 24.325 488.645 24.705 ;
        RECT 492.265 24.685 492.645 24.705 ;
        RECT 489.800 24.365 492.710 24.685 ;
        RECT 492.265 24.325 492.645 24.365 ;
        RECT 496.895 24.185 497.275 24.565 ;
        RECT 499.300 24.200 501.080 24.490 ;
        RECT 502.555 24.290 503.745 24.575 ;
        RECT 506.675 24.170 507.985 24.490 ;
        RECT 415.235 23.595 415.615 23.975 ;
        RECT 418.980 23.635 419.360 24.015 ;
        RECT 421.690 23.625 422.070 24.005 ;
        RECT 423.100 23.470 426.280 23.790 ;
        RECT 498.030 23.585 498.410 23.965 ;
        RECT 501.775 23.625 502.155 24.005 ;
        RECT 504.485 23.615 504.865 23.995 ;
        RECT 505.895 23.460 509.075 23.780 ;
        RECT 430.415 23.025 431.905 23.405 ;
        RECT 432.605 23.025 433.890 23.405 ;
        RECT 451.920 23.025 453.405 23.405 ;
        RECT 454.105 23.025 455.180 23.405 ;
        RECT 469.115 23.015 470.605 23.395 ;
        RECT 492.805 23.015 493.880 23.395 ;
        RECT 432.065 22.335 433.155 22.715 ;
        RECT 434.110 22.345 435.630 22.705 ;
        RECT 436.550 22.340 449.400 22.675 ;
        RECT 453.565 22.670 453.945 22.715 ;
        RECT 452.830 22.370 454.140 22.670 ;
        RECT 453.565 22.335 453.945 22.370 ;
        RECT 470.765 22.325 471.855 22.705 ;
        RECT 472.810 22.335 474.330 22.695 ;
        RECT 475.250 22.330 488.100 22.665 ;
        RECT 492.265 22.660 492.645 22.705 ;
        RECT 491.530 22.360 492.840 22.660 ;
        RECT 492.265 22.325 492.645 22.360 ;
        RECT 461.325 21.825 494.275 21.830 ;
        RECT 428.920 21.475 494.275 21.825 ;
        RECT 461.325 21.465 494.275 21.475 ;
        RECT 496.070 21.455 500.330 21.810 ;
        RECT 413.030 20.880 417.125 20.885 ;
        RECT 396.450 20.875 401.665 20.880 ;
        RECT 411.910 20.875 417.125 20.880 ;
        RECT 427.370 20.875 467.620 20.880 ;
        RECT 396.450 20.870 467.620 20.875 ;
        RECT 494.275 20.870 499.920 20.875 ;
        RECT 510.535 20.870 510.915 26.700 ;
        RECT 519.415 26.650 523.915 26.960 ;
        RECT 595.570 26.745 599.700 27.045 ;
        RECT 515.375 26.100 521.765 26.390 ;
        RECT 514.790 25.520 530.810 25.855 ;
        RECT 579.515 25.775 585.485 26.110 ;
        RECT 514.140 24.935 517.060 25.235 ;
        RECT 520.605 24.920 523.975 25.220 ;
        RECT 560.110 25.135 563.410 25.515 ;
        RECT 564.110 25.135 567.410 25.515 ;
        RECT 573.610 25.135 576.910 25.515 ;
        RECT 577.610 25.135 580.910 25.515 ;
        RECT 512.355 24.185 512.735 24.565 ;
        RECT 514.760 24.200 516.540 24.490 ;
        RECT 518.015 24.290 519.205 24.575 ;
        RECT 522.135 24.170 523.445 24.490 ;
        RECT 513.490 23.585 513.870 23.965 ;
        RECT 517.235 23.625 517.615 24.005 ;
        RECT 519.945 23.615 520.325 23.995 ;
        RECT 521.355 23.460 524.535 23.780 ;
        RECT 560.110 23.135 561.395 23.515 ;
        RECT 579.425 23.135 580.910 23.515 ;
        RECT 511.635 22.375 515.785 22.645 ;
        RECT 561.615 22.455 563.135 22.815 ;
        RECT 511.285 20.870 515.380 20.875 ;
        RECT 396.450 20.865 499.920 20.870 ;
        RECT 510.165 20.865 515.380 20.870 ;
        RECT 74.855 20.020 132.430 20.030 ;
        RECT 271.220 20.020 328.795 20.030 ;
        RECT 396.450 19.980 525.195 20.865 ;
        RECT 556.425 20.090 583.080 20.990 ;
        RECT 593.195 20.915 593.575 26.745 ;
        RECT 602.075 26.695 606.575 27.005 ;
        RECT 611.030 26.745 615.160 27.045 ;
        RECT 598.035 26.145 604.425 26.435 ;
        RECT 597.450 25.565 608.105 25.900 ;
        RECT 596.800 24.980 599.720 25.280 ;
        RECT 603.265 24.965 606.635 25.265 ;
        RECT 595.015 24.230 595.395 24.610 ;
        RECT 597.420 24.245 599.200 24.535 ;
        RECT 600.675 24.335 601.865 24.620 ;
        RECT 604.795 24.215 606.105 24.535 ;
        RECT 596.150 23.630 596.530 24.010 ;
        RECT 599.895 23.670 600.275 24.050 ;
        RECT 602.605 23.660 602.985 24.040 ;
        RECT 604.015 23.505 607.195 23.825 ;
        RECT 593.945 20.915 598.040 20.920 ;
        RECT 608.655 20.915 609.035 26.745 ;
        RECT 617.535 26.695 622.035 27.005 ;
        RECT 709.285 26.735 713.415 27.035 ;
        RECT 624.765 26.525 660.675 26.535 ;
        RECT 613.495 26.145 619.885 26.435 ;
        RECT 624.765 26.265 692.070 26.525 ;
        RECT 660.325 26.255 692.070 26.265 ;
        RECT 696.290 26.135 702.680 26.425 ;
        RECT 612.910 25.565 623.415 25.900 ;
        RECT 648.385 25.700 658.935 26.035 ;
        RECT 695.705 25.555 706.185 25.890 ;
        RECT 612.260 24.980 615.180 25.280 ;
        RECT 618.725 24.965 622.095 25.265 ;
        RECT 626.975 25.060 628.280 25.440 ;
        RECT 628.980 25.060 632.280 25.440 ;
        RECT 632.980 25.060 636.280 25.440 ;
        RECT 636.980 25.060 638.340 25.440 ;
        RECT 640.315 25.060 641.780 25.440 ;
        RECT 642.480 25.060 645.780 25.440 ;
        RECT 646.480 25.060 649.780 25.440 ;
        RECT 650.480 25.060 651.660 25.440 ;
        RECT 665.675 25.050 666.980 25.430 ;
        RECT 671.680 25.050 674.980 25.430 ;
        RECT 675.680 25.050 677.040 25.430 ;
        RECT 679.015 25.050 680.480 25.430 ;
        RECT 681.180 25.050 684.480 25.430 ;
        RECT 689.180 25.050 690.360 25.430 ;
        RECT 628.440 24.715 628.820 24.750 ;
        RECT 610.475 24.230 610.855 24.610 ;
        RECT 612.880 24.245 614.660 24.535 ;
        RECT 616.135 24.335 617.325 24.620 ;
        RECT 620.255 24.215 621.565 24.535 ;
        RECT 628.175 24.405 631.185 24.715 ;
        RECT 628.440 24.370 628.820 24.405 ;
        RECT 632.440 24.370 633.530 24.750 ;
        RECT 636.440 24.745 636.820 24.750 ;
        RECT 633.960 24.380 636.825 24.745 ;
        RECT 641.940 24.725 642.320 24.750 ;
        RECT 641.925 24.405 644.070 24.725 ;
        RECT 636.440 24.370 636.820 24.380 ;
        RECT 641.940 24.370 642.320 24.405 ;
        RECT 644.985 24.370 646.320 24.750 ;
        RECT 649.940 24.730 650.320 24.750 ;
        RECT 647.475 24.410 650.385 24.730 ;
        RECT 667.140 24.705 667.520 24.740 ;
        RECT 649.940 24.370 650.320 24.410 ;
        RECT 666.875 24.395 669.885 24.705 ;
        RECT 667.140 24.360 667.520 24.395 ;
        RECT 671.140 24.360 672.230 24.740 ;
        RECT 675.140 24.735 675.520 24.740 ;
        RECT 672.660 24.370 675.525 24.735 ;
        RECT 680.640 24.715 681.020 24.740 ;
        RECT 680.625 24.395 682.770 24.715 ;
        RECT 675.140 24.360 675.520 24.370 ;
        RECT 680.640 24.360 681.020 24.395 ;
        RECT 683.685 24.360 685.020 24.740 ;
        RECT 688.640 24.720 689.020 24.740 ;
        RECT 686.175 24.400 689.085 24.720 ;
        RECT 688.640 24.360 689.020 24.400 ;
        RECT 693.270 24.220 693.650 24.600 ;
        RECT 695.675 24.235 697.455 24.525 ;
        RECT 698.930 24.325 700.120 24.610 ;
        RECT 703.050 24.205 704.360 24.525 ;
        RECT 611.610 23.630 611.990 24.010 ;
        RECT 615.355 23.670 615.735 24.050 ;
        RECT 618.065 23.660 618.445 24.040 ;
        RECT 619.475 23.505 622.655 23.825 ;
        RECT 694.405 23.620 694.785 24.000 ;
        RECT 698.150 23.660 698.530 24.040 ;
        RECT 700.860 23.650 701.240 24.030 ;
        RECT 702.270 23.495 705.450 23.815 ;
        RECT 626.790 23.060 628.280 23.440 ;
        RECT 628.980 23.060 630.265 23.440 ;
        RECT 648.295 23.060 649.780 23.440 ;
        RECT 650.480 23.060 651.555 23.440 ;
        RECT 665.490 23.050 666.980 23.430 ;
        RECT 689.180 23.050 690.255 23.430 ;
        RECT 628.440 22.370 629.530 22.750 ;
        RECT 630.485 22.380 632.005 22.740 ;
        RECT 632.925 22.375 645.775 22.710 ;
        RECT 649.940 22.705 650.320 22.750 ;
        RECT 649.205 22.405 650.515 22.705 ;
        RECT 649.940 22.370 650.320 22.405 ;
        RECT 667.140 22.360 668.230 22.740 ;
        RECT 669.185 22.370 670.705 22.730 ;
        RECT 671.625 22.365 684.475 22.700 ;
        RECT 688.640 22.695 689.020 22.740 ;
        RECT 687.905 22.395 689.215 22.695 ;
        RECT 688.640 22.360 689.020 22.395 ;
        RECT 657.700 21.860 690.650 21.865 ;
        RECT 625.295 21.510 690.650 21.860 ;
        RECT 657.700 21.500 690.650 21.510 ;
        RECT 692.445 21.490 696.705 21.845 ;
        RECT 609.405 20.915 613.500 20.920 ;
        RECT 592.825 20.910 598.040 20.915 ;
        RECT 608.285 20.910 613.500 20.915 ;
        RECT 623.745 20.910 663.995 20.915 ;
        RECT 592.825 20.905 663.995 20.910 ;
        RECT 690.650 20.905 696.295 20.910 ;
        RECT 706.910 20.905 707.290 26.735 ;
        RECT 715.790 26.685 720.290 26.995 ;
        RECT 791.910 26.745 796.040 27.045 ;
        RECT 711.750 26.135 718.140 26.425 ;
        RECT 711.165 25.555 727.185 25.890 ;
        RECT 775.880 25.780 781.850 26.115 ;
        RECT 710.515 24.970 713.435 25.270 ;
        RECT 716.980 24.955 720.350 25.255 ;
        RECT 756.475 25.140 759.775 25.520 ;
        RECT 760.475 25.140 763.775 25.520 ;
        RECT 769.975 25.140 773.275 25.520 ;
        RECT 773.975 25.140 777.275 25.520 ;
        RECT 708.730 24.220 709.110 24.600 ;
        RECT 711.135 24.235 712.915 24.525 ;
        RECT 714.390 24.325 715.580 24.610 ;
        RECT 718.510 24.205 719.820 24.525 ;
        RECT 709.865 23.620 710.245 24.000 ;
        RECT 713.610 23.660 713.990 24.040 ;
        RECT 716.320 23.650 716.700 24.030 ;
        RECT 717.730 23.495 720.910 23.815 ;
        RECT 756.475 23.140 757.760 23.520 ;
        RECT 775.790 23.140 777.275 23.520 ;
        RECT 708.010 22.410 712.160 22.680 ;
        RECT 757.980 22.460 759.500 22.820 ;
        RECT 707.660 20.905 711.755 20.910 ;
        RECT 592.825 20.900 696.295 20.905 ;
        RECT 706.540 20.900 711.755 20.905 ;
        RECT 592.825 20.015 721.570 20.900 ;
        RECT 752.790 20.095 779.445 20.995 ;
        RECT 789.535 20.915 789.915 26.745 ;
        RECT 798.415 26.695 802.915 27.005 ;
        RECT 807.370 26.745 811.500 27.045 ;
        RECT 794.375 26.145 800.765 26.435 ;
        RECT 793.790 25.565 804.445 25.900 ;
        RECT 793.140 24.980 796.060 25.280 ;
        RECT 799.605 24.965 802.975 25.265 ;
        RECT 791.355 24.230 791.735 24.610 ;
        RECT 793.760 24.245 795.540 24.535 ;
        RECT 797.015 24.335 798.205 24.620 ;
        RECT 801.135 24.215 802.445 24.535 ;
        RECT 792.490 23.630 792.870 24.010 ;
        RECT 796.235 23.670 796.615 24.050 ;
        RECT 798.945 23.660 799.325 24.040 ;
        RECT 800.355 23.505 803.535 23.825 ;
        RECT 790.285 20.915 794.380 20.920 ;
        RECT 804.995 20.915 805.375 26.745 ;
        RECT 813.875 26.695 818.375 27.005 ;
        RECT 905.625 26.735 909.755 27.035 ;
        RECT 821.105 26.525 857.015 26.535 ;
        RECT 809.835 26.145 816.225 26.435 ;
        RECT 821.105 26.265 888.410 26.525 ;
        RECT 856.665 26.255 888.410 26.265 ;
        RECT 892.630 26.135 899.020 26.425 ;
        RECT 809.250 25.565 819.755 25.900 ;
        RECT 844.725 25.700 855.275 26.035 ;
        RECT 892.045 25.555 902.525 25.890 ;
        RECT 808.600 24.980 811.520 25.280 ;
        RECT 815.065 24.965 818.435 25.265 ;
        RECT 823.315 25.060 824.620 25.440 ;
        RECT 825.320 25.060 828.620 25.440 ;
        RECT 829.320 25.060 832.620 25.440 ;
        RECT 833.320 25.060 834.680 25.440 ;
        RECT 836.655 25.060 838.120 25.440 ;
        RECT 838.820 25.060 842.120 25.440 ;
        RECT 842.820 25.060 846.120 25.440 ;
        RECT 846.820 25.060 848.000 25.440 ;
        RECT 862.015 25.050 863.320 25.430 ;
        RECT 868.020 25.050 871.320 25.430 ;
        RECT 872.020 25.050 873.380 25.430 ;
        RECT 875.355 25.050 876.820 25.430 ;
        RECT 877.520 25.050 880.820 25.430 ;
        RECT 885.520 25.050 886.700 25.430 ;
        RECT 824.780 24.715 825.160 24.750 ;
        RECT 806.815 24.230 807.195 24.610 ;
        RECT 809.220 24.245 811.000 24.535 ;
        RECT 812.475 24.335 813.665 24.620 ;
        RECT 816.595 24.215 817.905 24.535 ;
        RECT 824.515 24.405 827.525 24.715 ;
        RECT 824.780 24.370 825.160 24.405 ;
        RECT 828.780 24.370 829.870 24.750 ;
        RECT 832.780 24.745 833.160 24.750 ;
        RECT 830.300 24.380 833.165 24.745 ;
        RECT 838.280 24.725 838.660 24.750 ;
        RECT 838.265 24.405 840.410 24.725 ;
        RECT 832.780 24.370 833.160 24.380 ;
        RECT 838.280 24.370 838.660 24.405 ;
        RECT 841.325 24.370 842.660 24.750 ;
        RECT 846.280 24.730 846.660 24.750 ;
        RECT 843.815 24.410 846.725 24.730 ;
        RECT 863.480 24.705 863.860 24.740 ;
        RECT 846.280 24.370 846.660 24.410 ;
        RECT 863.215 24.395 866.225 24.705 ;
        RECT 863.480 24.360 863.860 24.395 ;
        RECT 867.480 24.360 868.570 24.740 ;
        RECT 871.480 24.735 871.860 24.740 ;
        RECT 869.000 24.370 871.865 24.735 ;
        RECT 876.980 24.715 877.360 24.740 ;
        RECT 876.965 24.395 879.110 24.715 ;
        RECT 871.480 24.360 871.860 24.370 ;
        RECT 876.980 24.360 877.360 24.395 ;
        RECT 880.025 24.360 881.360 24.740 ;
        RECT 884.980 24.720 885.360 24.740 ;
        RECT 882.515 24.400 885.425 24.720 ;
        RECT 884.980 24.360 885.360 24.400 ;
        RECT 889.610 24.220 889.990 24.600 ;
        RECT 892.015 24.235 893.795 24.525 ;
        RECT 895.270 24.325 896.460 24.610 ;
        RECT 899.390 24.205 900.700 24.525 ;
        RECT 807.950 23.630 808.330 24.010 ;
        RECT 811.695 23.670 812.075 24.050 ;
        RECT 814.405 23.660 814.785 24.040 ;
        RECT 815.815 23.505 818.995 23.825 ;
        RECT 890.745 23.620 891.125 24.000 ;
        RECT 894.490 23.660 894.870 24.040 ;
        RECT 897.200 23.650 897.580 24.030 ;
        RECT 898.610 23.495 901.790 23.815 ;
        RECT 823.130 23.060 824.620 23.440 ;
        RECT 825.320 23.060 826.605 23.440 ;
        RECT 844.635 23.060 846.120 23.440 ;
        RECT 846.820 23.060 847.895 23.440 ;
        RECT 861.830 23.050 863.320 23.430 ;
        RECT 885.520 23.050 886.595 23.430 ;
        RECT 824.780 22.370 825.870 22.750 ;
        RECT 826.825 22.380 828.345 22.740 ;
        RECT 829.265 22.375 842.115 22.710 ;
        RECT 846.280 22.705 846.660 22.750 ;
        RECT 845.545 22.405 846.855 22.705 ;
        RECT 846.280 22.370 846.660 22.405 ;
        RECT 863.480 22.360 864.570 22.740 ;
        RECT 865.525 22.370 867.045 22.730 ;
        RECT 867.965 22.365 880.815 22.700 ;
        RECT 884.980 22.695 885.360 22.740 ;
        RECT 884.245 22.395 885.555 22.695 ;
        RECT 884.980 22.360 885.360 22.395 ;
        RECT 854.040 21.860 886.990 21.865 ;
        RECT 821.635 21.510 886.990 21.860 ;
        RECT 854.040 21.500 886.990 21.510 ;
        RECT 888.785 21.490 893.045 21.845 ;
        RECT 805.745 20.915 809.840 20.920 ;
        RECT 789.165 20.910 794.380 20.915 ;
        RECT 804.625 20.910 809.840 20.915 ;
        RECT 820.085 20.910 860.335 20.915 ;
        RECT 789.165 20.905 860.335 20.910 ;
        RECT 886.990 20.905 892.635 20.910 ;
        RECT 903.250 20.905 903.630 26.735 ;
        RECT 912.130 26.685 916.630 26.995 ;
        RECT 988.250 26.745 992.380 27.045 ;
        RECT 908.090 26.135 914.480 26.425 ;
        RECT 907.505 25.555 923.525 25.890 ;
        RECT 972.265 25.765 978.235 26.100 ;
        RECT 906.855 24.970 909.775 25.270 ;
        RECT 913.320 24.955 916.690 25.255 ;
        RECT 952.860 25.125 956.160 25.505 ;
        RECT 956.860 25.125 960.160 25.505 ;
        RECT 966.360 25.125 969.660 25.505 ;
        RECT 970.360 25.125 973.660 25.505 ;
        RECT 905.070 24.220 905.450 24.600 ;
        RECT 907.475 24.235 909.255 24.525 ;
        RECT 910.730 24.325 911.920 24.610 ;
        RECT 914.850 24.205 916.160 24.525 ;
        RECT 906.205 23.620 906.585 24.000 ;
        RECT 909.950 23.660 910.330 24.040 ;
        RECT 912.660 23.650 913.040 24.030 ;
        RECT 914.070 23.495 917.250 23.815 ;
        RECT 952.860 23.125 954.145 23.505 ;
        RECT 972.175 23.125 973.660 23.505 ;
        RECT 904.350 22.410 908.500 22.680 ;
        RECT 954.365 22.445 955.885 22.805 ;
        RECT 904.000 20.905 908.095 20.910 ;
        RECT 789.165 20.900 892.635 20.905 ;
        RECT 902.880 20.900 908.095 20.905 ;
        RECT 789.165 20.015 917.910 20.900 ;
        RECT 949.175 20.080 975.830 20.980 ;
        RECT 985.875 20.915 986.255 26.745 ;
        RECT 994.755 26.695 999.255 27.005 ;
        RECT 1003.710 26.745 1007.840 27.045 ;
        RECT 990.715 26.145 997.105 26.435 ;
        RECT 990.130 25.565 1000.785 25.900 ;
        RECT 989.480 24.980 992.400 25.280 ;
        RECT 995.945 24.965 999.315 25.265 ;
        RECT 987.695 24.230 988.075 24.610 ;
        RECT 990.100 24.245 991.880 24.535 ;
        RECT 993.355 24.335 994.545 24.620 ;
        RECT 997.475 24.215 998.785 24.535 ;
        RECT 988.830 23.630 989.210 24.010 ;
        RECT 992.575 23.670 992.955 24.050 ;
        RECT 995.285 23.660 995.665 24.040 ;
        RECT 996.695 23.505 999.875 23.825 ;
        RECT 986.625 20.915 990.720 20.920 ;
        RECT 1001.335 20.915 1001.715 26.745 ;
        RECT 1010.215 26.695 1014.715 27.005 ;
        RECT 1101.965 26.735 1106.095 27.035 ;
        RECT 1017.445 26.525 1053.355 26.535 ;
        RECT 1006.175 26.145 1012.565 26.435 ;
        RECT 1017.445 26.265 1084.750 26.525 ;
        RECT 1053.005 26.255 1084.750 26.265 ;
        RECT 1088.970 26.135 1095.360 26.425 ;
        RECT 1005.590 25.565 1016.095 25.900 ;
        RECT 1041.065 25.700 1051.615 26.035 ;
        RECT 1088.385 25.555 1098.865 25.890 ;
        RECT 1004.940 24.980 1007.860 25.280 ;
        RECT 1011.405 24.965 1014.775 25.265 ;
        RECT 1019.655 25.060 1020.960 25.440 ;
        RECT 1021.660 25.060 1024.960 25.440 ;
        RECT 1025.660 25.060 1028.960 25.440 ;
        RECT 1029.660 25.060 1031.020 25.440 ;
        RECT 1032.995 25.060 1034.460 25.440 ;
        RECT 1035.160 25.060 1038.460 25.440 ;
        RECT 1039.160 25.060 1042.460 25.440 ;
        RECT 1043.160 25.060 1044.340 25.440 ;
        RECT 1058.355 25.050 1059.660 25.430 ;
        RECT 1064.360 25.050 1067.660 25.430 ;
        RECT 1068.360 25.050 1069.720 25.430 ;
        RECT 1071.695 25.050 1073.160 25.430 ;
        RECT 1073.860 25.050 1077.160 25.430 ;
        RECT 1081.860 25.050 1083.040 25.430 ;
        RECT 1021.120 24.715 1021.500 24.750 ;
        RECT 1003.155 24.230 1003.535 24.610 ;
        RECT 1005.560 24.245 1007.340 24.535 ;
        RECT 1008.815 24.335 1010.005 24.620 ;
        RECT 1012.935 24.215 1014.245 24.535 ;
        RECT 1020.855 24.405 1023.865 24.715 ;
        RECT 1021.120 24.370 1021.500 24.405 ;
        RECT 1025.120 24.370 1026.210 24.750 ;
        RECT 1029.120 24.745 1029.500 24.750 ;
        RECT 1026.640 24.380 1029.505 24.745 ;
        RECT 1034.620 24.725 1035.000 24.750 ;
        RECT 1034.605 24.405 1036.750 24.725 ;
        RECT 1029.120 24.370 1029.500 24.380 ;
        RECT 1034.620 24.370 1035.000 24.405 ;
        RECT 1037.665 24.370 1039.000 24.750 ;
        RECT 1042.620 24.730 1043.000 24.750 ;
        RECT 1040.155 24.410 1043.065 24.730 ;
        RECT 1059.820 24.705 1060.200 24.740 ;
        RECT 1042.620 24.370 1043.000 24.410 ;
        RECT 1059.555 24.395 1062.565 24.705 ;
        RECT 1059.820 24.360 1060.200 24.395 ;
        RECT 1063.820 24.360 1064.910 24.740 ;
        RECT 1067.820 24.735 1068.200 24.740 ;
        RECT 1065.340 24.370 1068.205 24.735 ;
        RECT 1073.320 24.715 1073.700 24.740 ;
        RECT 1073.305 24.395 1075.450 24.715 ;
        RECT 1067.820 24.360 1068.200 24.370 ;
        RECT 1073.320 24.360 1073.700 24.395 ;
        RECT 1076.365 24.360 1077.700 24.740 ;
        RECT 1081.320 24.720 1081.700 24.740 ;
        RECT 1078.855 24.400 1081.765 24.720 ;
        RECT 1081.320 24.360 1081.700 24.400 ;
        RECT 1085.950 24.220 1086.330 24.600 ;
        RECT 1088.355 24.235 1090.135 24.525 ;
        RECT 1091.610 24.325 1092.800 24.610 ;
        RECT 1095.730 24.205 1097.040 24.525 ;
        RECT 1004.290 23.630 1004.670 24.010 ;
        RECT 1008.035 23.670 1008.415 24.050 ;
        RECT 1010.745 23.660 1011.125 24.040 ;
        RECT 1012.155 23.505 1015.335 23.825 ;
        RECT 1087.085 23.620 1087.465 24.000 ;
        RECT 1090.830 23.660 1091.210 24.040 ;
        RECT 1093.540 23.650 1093.920 24.030 ;
        RECT 1094.950 23.495 1098.130 23.815 ;
        RECT 1019.470 23.060 1020.960 23.440 ;
        RECT 1021.660 23.060 1022.945 23.440 ;
        RECT 1040.975 23.060 1042.460 23.440 ;
        RECT 1043.160 23.060 1044.235 23.440 ;
        RECT 1058.170 23.050 1059.660 23.430 ;
        RECT 1081.860 23.050 1082.935 23.430 ;
        RECT 1021.120 22.370 1022.210 22.750 ;
        RECT 1023.165 22.380 1024.685 22.740 ;
        RECT 1025.605 22.375 1038.455 22.710 ;
        RECT 1042.620 22.705 1043.000 22.750 ;
        RECT 1041.885 22.405 1043.195 22.705 ;
        RECT 1042.620 22.370 1043.000 22.405 ;
        RECT 1059.820 22.360 1060.910 22.740 ;
        RECT 1061.865 22.370 1063.385 22.730 ;
        RECT 1064.305 22.365 1077.155 22.700 ;
        RECT 1081.320 22.695 1081.700 22.740 ;
        RECT 1080.585 22.395 1081.895 22.695 ;
        RECT 1081.320 22.360 1081.700 22.395 ;
        RECT 1050.380 21.860 1083.330 21.865 ;
        RECT 1017.975 21.510 1083.330 21.860 ;
        RECT 1050.380 21.500 1083.330 21.510 ;
        RECT 1085.125 21.490 1089.385 21.845 ;
        RECT 1002.085 20.915 1006.180 20.920 ;
        RECT 985.505 20.910 990.720 20.915 ;
        RECT 1000.965 20.910 1006.180 20.915 ;
        RECT 1016.425 20.910 1056.675 20.915 ;
        RECT 985.505 20.905 1056.675 20.910 ;
        RECT 1083.330 20.905 1088.975 20.910 ;
        RECT 1099.590 20.905 1099.970 26.735 ;
        RECT 1108.470 26.685 1112.970 26.995 ;
        RECT 1184.590 26.745 1188.720 27.045 ;
        RECT 1104.430 26.135 1110.820 26.425 ;
        RECT 1103.845 25.555 1119.865 25.890 ;
        RECT 1168.590 25.770 1174.560 26.105 ;
        RECT 1103.195 24.970 1106.115 25.270 ;
        RECT 1109.660 24.955 1113.030 25.255 ;
        RECT 1149.185 25.130 1152.485 25.510 ;
        RECT 1153.185 25.130 1156.485 25.510 ;
        RECT 1162.685 25.130 1165.985 25.510 ;
        RECT 1166.685 25.130 1169.985 25.510 ;
        RECT 1101.410 24.220 1101.790 24.600 ;
        RECT 1103.815 24.235 1105.595 24.525 ;
        RECT 1107.070 24.325 1108.260 24.610 ;
        RECT 1111.190 24.205 1112.500 24.525 ;
        RECT 1102.545 23.620 1102.925 24.000 ;
        RECT 1106.290 23.660 1106.670 24.040 ;
        RECT 1109.000 23.650 1109.380 24.030 ;
        RECT 1110.410 23.495 1113.590 23.815 ;
        RECT 1149.185 23.130 1150.470 23.510 ;
        RECT 1168.500 23.130 1169.985 23.510 ;
        RECT 1100.690 22.410 1104.840 22.680 ;
        RECT 1150.690 22.450 1152.210 22.810 ;
        RECT 1100.340 20.905 1104.435 20.910 ;
        RECT 985.505 20.900 1088.975 20.905 ;
        RECT 1099.220 20.900 1104.435 20.905 ;
        RECT 985.505 20.015 1114.250 20.900 ;
        RECT 1145.500 20.085 1172.155 20.985 ;
        RECT 1182.215 20.915 1182.595 26.745 ;
        RECT 1191.095 26.695 1195.595 27.005 ;
        RECT 1200.050 26.745 1204.180 27.045 ;
        RECT 1187.055 26.145 1193.445 26.435 ;
        RECT 1186.470 25.565 1197.125 25.900 ;
        RECT 1185.820 24.980 1188.740 25.280 ;
        RECT 1192.285 24.965 1195.655 25.265 ;
        RECT 1184.035 24.230 1184.415 24.610 ;
        RECT 1186.440 24.245 1188.220 24.535 ;
        RECT 1189.695 24.335 1190.885 24.620 ;
        RECT 1193.815 24.215 1195.125 24.535 ;
        RECT 1185.170 23.630 1185.550 24.010 ;
        RECT 1188.915 23.670 1189.295 24.050 ;
        RECT 1191.625 23.660 1192.005 24.040 ;
        RECT 1193.035 23.505 1196.215 23.825 ;
        RECT 1182.965 20.915 1187.060 20.920 ;
        RECT 1197.675 20.915 1198.055 26.745 ;
        RECT 1206.555 26.695 1211.055 27.005 ;
        RECT 1282.845 26.735 1286.975 27.035 ;
        RECT 1289.350 26.685 1293.850 26.995 ;
        RECT 1298.305 26.735 1302.435 27.035 ;
        RECT 1213.785 26.525 1249.695 26.535 ;
        RECT 1202.515 26.145 1208.905 26.435 ;
        RECT 1213.785 26.265 1281.090 26.525 ;
        RECT 1249.345 26.255 1281.090 26.265 ;
        RECT 1285.310 26.135 1291.700 26.425 ;
        RECT 1201.930 25.565 1212.435 25.900 ;
        RECT 1237.405 25.700 1247.955 26.035 ;
        RECT 1276.105 25.690 1280.050 26.025 ;
        RECT 1284.725 25.555 1295.205 25.890 ;
        RECT 1201.280 24.980 1204.200 25.280 ;
        RECT 1207.745 24.965 1211.115 25.265 ;
        RECT 1215.995 25.060 1217.300 25.440 ;
        RECT 1218.000 25.060 1221.300 25.440 ;
        RECT 1222.000 25.060 1225.300 25.440 ;
        RECT 1226.000 25.060 1227.360 25.440 ;
        RECT 1229.335 25.060 1230.800 25.440 ;
        RECT 1231.500 25.060 1234.800 25.440 ;
        RECT 1235.500 25.060 1238.800 25.440 ;
        RECT 1239.500 25.060 1240.680 25.440 ;
        RECT 1254.695 25.050 1256.000 25.430 ;
        RECT 1256.700 25.050 1260.000 25.430 ;
        RECT 1260.700 25.050 1264.000 25.430 ;
        RECT 1264.700 25.050 1266.060 25.430 ;
        RECT 1268.035 25.050 1269.500 25.430 ;
        RECT 1270.200 25.050 1273.500 25.430 ;
        RECT 1274.200 25.050 1277.500 25.430 ;
        RECT 1278.200 25.050 1279.380 25.430 ;
        RECT 1284.075 24.970 1286.995 25.270 ;
        RECT 1290.540 24.955 1293.910 25.255 ;
        RECT 1217.460 24.715 1217.840 24.750 ;
        RECT 1199.495 24.230 1199.875 24.610 ;
        RECT 1201.900 24.245 1203.680 24.535 ;
        RECT 1205.155 24.335 1206.345 24.620 ;
        RECT 1209.275 24.215 1210.585 24.535 ;
        RECT 1217.195 24.405 1220.205 24.715 ;
        RECT 1217.460 24.370 1217.840 24.405 ;
        RECT 1221.460 24.370 1222.550 24.750 ;
        RECT 1225.460 24.745 1225.840 24.750 ;
        RECT 1222.980 24.380 1225.845 24.745 ;
        RECT 1230.960 24.725 1231.340 24.750 ;
        RECT 1230.945 24.405 1233.090 24.725 ;
        RECT 1225.460 24.370 1225.840 24.380 ;
        RECT 1230.960 24.370 1231.340 24.405 ;
        RECT 1234.005 24.370 1235.340 24.750 ;
        RECT 1238.960 24.730 1239.340 24.750 ;
        RECT 1236.495 24.410 1239.405 24.730 ;
        RECT 1256.160 24.705 1256.540 24.740 ;
        RECT 1238.960 24.370 1239.340 24.410 ;
        RECT 1255.895 24.395 1258.905 24.705 ;
        RECT 1256.160 24.360 1256.540 24.395 ;
        RECT 1260.160 24.360 1261.250 24.740 ;
        RECT 1264.160 24.735 1264.540 24.740 ;
        RECT 1261.680 24.370 1264.545 24.735 ;
        RECT 1269.660 24.715 1270.040 24.740 ;
        RECT 1269.645 24.395 1271.790 24.715 ;
        RECT 1264.160 24.360 1264.540 24.370 ;
        RECT 1269.660 24.360 1270.040 24.395 ;
        RECT 1272.705 24.360 1274.040 24.740 ;
        RECT 1277.660 24.720 1278.040 24.740 ;
        RECT 1275.195 24.400 1278.105 24.720 ;
        RECT 1277.660 24.360 1278.040 24.400 ;
        RECT 1282.290 24.220 1282.670 24.600 ;
        RECT 1284.695 24.235 1286.475 24.525 ;
        RECT 1287.950 24.325 1289.140 24.610 ;
        RECT 1292.070 24.205 1293.380 24.525 ;
        RECT 1200.630 23.630 1201.010 24.010 ;
        RECT 1204.375 23.670 1204.755 24.050 ;
        RECT 1207.085 23.660 1207.465 24.040 ;
        RECT 1208.495 23.505 1211.675 23.825 ;
        RECT 1283.425 23.620 1283.805 24.000 ;
        RECT 1287.170 23.660 1287.550 24.040 ;
        RECT 1289.880 23.650 1290.260 24.030 ;
        RECT 1291.290 23.495 1294.470 23.815 ;
        RECT 1215.810 23.060 1217.300 23.440 ;
        RECT 1218.000 23.060 1219.285 23.440 ;
        RECT 1237.315 23.060 1238.800 23.440 ;
        RECT 1239.500 23.060 1240.575 23.440 ;
        RECT 1254.510 23.050 1256.000 23.430 ;
        RECT 1256.700 23.050 1257.985 23.430 ;
        RECT 1276.015 23.050 1277.500 23.430 ;
        RECT 1278.200 23.050 1279.275 23.430 ;
        RECT 1217.460 22.370 1218.550 22.750 ;
        RECT 1219.505 22.380 1221.025 22.740 ;
        RECT 1221.945 22.375 1234.795 22.710 ;
        RECT 1238.960 22.705 1239.340 22.750 ;
        RECT 1238.225 22.405 1239.535 22.705 ;
        RECT 1238.960 22.370 1239.340 22.405 ;
        RECT 1256.160 22.360 1257.250 22.740 ;
        RECT 1258.205 22.370 1259.725 22.730 ;
        RECT 1260.645 22.365 1273.495 22.700 ;
        RECT 1277.660 22.695 1278.040 22.740 ;
        RECT 1276.925 22.395 1278.235 22.695 ;
        RECT 1277.660 22.360 1278.040 22.395 ;
        RECT 1246.720 21.860 1279.670 21.865 ;
        RECT 1214.315 21.510 1279.670 21.860 ;
        RECT 1246.720 21.500 1279.670 21.510 ;
        RECT 1281.465 21.490 1285.725 21.845 ;
        RECT 1198.425 20.915 1202.520 20.920 ;
        RECT 1181.845 20.910 1187.060 20.915 ;
        RECT 1197.305 20.910 1202.520 20.915 ;
        RECT 1212.765 20.910 1253.015 20.915 ;
        RECT 1181.845 20.905 1253.015 20.910 ;
        RECT 1279.670 20.905 1285.315 20.910 ;
        RECT 1295.930 20.905 1296.310 26.735 ;
        RECT 1304.810 26.685 1309.310 26.995 ;
        RECT 1300.770 26.135 1307.160 26.425 ;
        RECT 1299.535 24.970 1302.455 25.270 ;
        RECT 1306.000 24.955 1309.370 25.255 ;
        RECT 1297.750 24.220 1298.130 24.600 ;
        RECT 1303.410 24.325 1304.600 24.610 ;
        RECT 1302.630 23.660 1303.010 24.040 ;
        RECT 1306.750 23.495 1309.930 23.815 ;
        RECT 1297.030 22.410 1301.180 22.680 ;
        RECT 1296.680 20.905 1300.775 20.910 ;
        RECT 1181.845 20.900 1285.315 20.905 ;
        RECT 1295.560 20.900 1300.775 20.905 ;
        RECT 1181.845 20.015 1310.590 20.900 ;
        RECT 663.995 20.005 721.570 20.015 ;
        RECT 860.335 20.005 917.910 20.015 ;
        RECT 1056.675 20.005 1114.250 20.015 ;
        RECT 1253.015 20.005 1310.590 20.015 ;
        RECT 467.620 19.970 525.195 19.980 ;
        RECT 79.265 10.855 79.645 11.235 ;
        RECT 86.165 10.845 86.545 11.225 ;
        RECT 275.630 10.855 276.010 11.235 ;
        RECT 282.530 10.845 282.910 11.225 ;
        RECT 472.030 10.805 472.410 11.185 ;
        RECT 478.930 10.795 479.310 11.175 ;
        RECT 668.405 10.840 668.785 11.220 ;
        RECT 675.305 10.830 675.685 11.210 ;
        RECT 864.745 10.840 865.125 11.220 ;
        RECT 871.645 10.830 872.025 11.210 ;
        RECT 1061.085 10.840 1061.465 11.220 ;
        RECT 1067.985 10.830 1068.365 11.210 ;
        RECT 76.590 10.430 78.330 10.720 ;
        RECT 83.090 10.375 85.680 10.725 ;
        RECT 272.955 10.430 274.695 10.720 ;
        RECT 279.455 10.375 282.045 10.725 ;
        RECT 469.355 10.380 471.095 10.670 ;
        RECT 475.855 10.325 478.445 10.675 ;
        RECT 665.730 10.415 667.470 10.705 ;
        RECT 672.230 10.360 674.820 10.710 ;
        RECT 862.070 10.415 863.810 10.705 ;
        RECT 868.570 10.360 871.160 10.710 ;
        RECT 1058.410 10.415 1060.150 10.705 ;
        RECT 1064.910 10.360 1067.500 10.710 ;
        RECT 71.025 9.670 88.350 9.970 ;
        RECT 267.390 9.670 284.715 9.970 ;
        RECT 463.790 9.620 481.115 9.920 ;
        RECT 660.165 9.655 677.490 9.955 ;
        RECT 856.505 9.655 873.830 9.955 ;
        RECT 1052.845 9.655 1070.170 9.955 ;
        RECT 1249.185 9.655 1266.510 9.955 ;
        RECT 70.785 8.925 88.350 9.225 ;
        RECT 267.150 8.925 284.715 9.225 ;
        RECT 463.550 8.875 481.115 9.175 ;
        RECT 659.925 8.910 677.490 9.210 ;
        RECT 856.265 8.910 873.830 9.210 ;
        RECT 1052.605 8.910 1070.170 9.210 ;
        RECT 1248.945 8.910 1266.510 9.210 ;
        RECT 85.275 7.910 88.350 8.185 ;
        RECT 281.640 7.910 284.715 8.185 ;
        RECT 478.040 7.860 481.115 8.135 ;
        RECT 674.415 7.895 677.490 8.170 ;
        RECT 870.755 7.895 873.830 8.170 ;
        RECT 1067.095 7.895 1070.170 8.170 ;
        RECT 76.065 7.015 80.195 7.315 ;
        RECT 82.570 6.965 87.070 7.275 ;
        RECT 272.430 7.015 276.560 7.315 ;
        RECT 278.935 6.965 283.435 7.275 ;
        RECT 468.830 6.965 472.960 7.265 ;
        RECT 475.335 6.915 479.835 7.225 ;
        RECT 665.205 7.000 669.335 7.300 ;
        RECT 671.710 6.950 676.210 7.260 ;
        RECT 861.545 7.000 865.675 7.300 ;
        RECT 868.050 6.950 872.550 7.260 ;
        RECT 1057.885 7.000 1062.015 7.300 ;
        RECT 1064.390 6.950 1068.890 7.260 ;
        RECT 1254.225 7.000 1258.355 7.300 ;
        RECT 1260.730 6.950 1265.230 7.260 ;
        RECT 77.945 5.835 88.350 6.170 ;
        RECT 274.310 5.835 284.715 6.170 ;
        RECT 470.710 5.785 481.115 6.120 ;
        RECT 667.085 5.820 677.490 6.155 ;
        RECT 863.425 5.820 873.830 6.155 ;
        RECT 1059.765 5.820 1070.170 6.155 ;
        RECT 77.295 5.250 80.215 5.550 ;
        RECT 83.760 5.235 87.130 5.535 ;
        RECT 273.660 5.250 276.580 5.550 ;
        RECT 280.125 5.235 283.495 5.535 ;
        RECT 470.060 5.200 472.980 5.500 ;
        RECT 476.525 5.185 479.895 5.485 ;
        RECT 666.435 5.235 669.355 5.535 ;
        RECT 672.900 5.220 676.270 5.520 ;
        RECT 862.775 5.235 865.695 5.535 ;
        RECT 869.240 5.220 872.610 5.520 ;
        RECT 1059.115 5.235 1062.035 5.535 ;
        RECT 1065.580 5.220 1068.950 5.520 ;
        RECT 1255.455 5.235 1258.375 5.535 ;
        RECT 1261.920 5.220 1265.290 5.520 ;
        RECT 77.915 4.515 79.695 4.805 ;
        RECT 85.290 4.485 86.600 4.805 ;
        RECT 274.280 4.515 276.060 4.805 ;
        RECT 281.655 4.485 282.965 4.805 ;
        RECT 470.680 4.465 472.460 4.755 ;
        RECT 478.055 4.435 479.365 4.755 ;
        RECT 667.055 4.500 668.835 4.790 ;
        RECT 674.430 4.470 675.740 4.790 ;
        RECT 863.395 4.500 865.175 4.790 ;
        RECT 870.770 4.470 872.080 4.790 ;
        RECT 1059.735 4.500 1061.515 4.790 ;
        RECT 1067.110 4.470 1068.420 4.790 ;
        RECT 76.645 3.900 77.025 4.280 ;
        RECT 83.100 3.930 83.480 4.310 ;
        RECT 273.010 3.900 273.390 4.280 ;
        RECT 279.465 3.930 279.845 4.310 ;
        RECT 469.410 3.850 469.790 4.230 ;
        RECT 475.865 3.880 476.245 4.260 ;
        RECT 665.785 3.885 666.165 4.265 ;
        RECT 672.240 3.915 672.620 4.295 ;
        RECT 862.125 3.885 862.505 4.265 ;
        RECT 868.580 3.915 868.960 4.295 ;
        RECT 1058.465 3.885 1058.845 4.265 ;
        RECT 1064.920 3.915 1065.300 4.295 ;
      LAYER Metal2 ;
        RECT -24.090 190.685 -23.690 193.735 ;
        RECT -19.170 190.595 -18.760 193.690 ;
        RECT -14.590 190.570 -14.180 193.665 ;
        RECT -26.255 178.490 -25.910 180.950 ;
        RECT -78.160 160.605 -77.845 171.655 ;
        RECT -74.325 170.950 -73.925 174.000 ;
        RECT -69.405 170.860 -68.995 173.955 ;
        RECT -64.825 170.835 -64.415 173.930 ;
        RECT -76.490 158.755 -76.145 161.215 ;
        RECT -59.375 161.090 -59.060 171.775 ;
        RECT -55.685 163.885 -55.270 166.700 ;
        RECT -54.945 165.470 -54.560 167.365 ;
        RECT -27.835 160.685 -27.520 171.735 ;
        RECT -24.000 171.030 -23.600 174.080 ;
        RECT -19.080 170.940 -18.670 174.035 ;
        RECT -14.500 170.915 -14.090 174.010 ;
        RECT -26.165 158.835 -25.820 161.295 ;
        RECT -9.050 161.170 -8.735 171.855 ;
        RECT -3.865 163.960 -3.415 168.120 ;
        RECT 5.335 167.685 5.715 168.065 ;
        RECT -2.165 166.940 -1.640 167.380 ;
        RECT 5.325 166.935 5.705 167.315 ;
        RECT 5.370 166.250 5.750 166.630 ;
        RECT 5.335 165.580 5.715 165.960 ;
        RECT 6.050 162.505 6.350 169.545 ;
        RECT 7.170 161.900 7.470 168.830 ;
        RECT 7.825 163.260 8.125 167.320 ;
        RECT 8.480 162.500 8.780 168.850 ;
        RECT 9.075 164.375 9.395 169.535 ;
        RECT 9.795 162.530 10.090 169.355 ;
        RECT 10.925 161.990 11.225 168.800 ;
        RECT 11.715 162.585 12.025 168.775 ;
        RECT 12.510 162.515 12.810 169.345 ;
        RECT 13.635 161.900 13.935 168.840 ;
        RECT 14.315 163.245 14.595 167.335 ;
        RECT 15.085 161.775 15.365 164.810 ;
        RECT 15.845 162.475 16.150 168.835 ;
        RECT 16.695 162.475 16.995 169.295 ;
        RECT 17.835 161.730 18.135 168.885 ;
        RECT 18.500 167.685 18.880 168.065 ;
        RECT 20.770 167.685 21.150 168.090 ;
        RECT 18.505 166.935 18.885 167.315 ;
        RECT 20.775 166.935 21.155 167.340 ;
        RECT 18.505 165.920 18.885 166.300 ;
        RECT 18.720 161.210 19.100 164.230 ;
        RECT 22.630 161.900 22.930 168.830 ;
        RECT 23.285 163.260 23.585 167.320 ;
        RECT 23.940 162.500 24.240 168.850 ;
        RECT 25.255 162.530 25.550 169.355 ;
        RECT 29.095 161.900 29.395 168.840 ;
        RECT 29.775 163.245 30.055 167.335 ;
        RECT 31.305 162.475 31.625 168.835 ;
        RECT 32.155 162.475 32.455 169.295 ;
        RECT 34.235 167.685 34.595 169.515 ;
        RECT 33.930 163.875 34.310 164.255 ;
        RECT 34.635 159.760 34.995 166.320 ;
        RECT 35.775 164.510 36.100 166.375 ;
        RECT 36.415 166.165 36.830 169.515 ;
        RECT 36.440 161.165 36.900 165.850 ;
        RECT 37.225 163.710 37.675 172.530 ;
        RECT 38.085 161.335 38.440 171.640 ;
        RECT 38.750 166.940 39.095 167.995 ;
        RECT 39.410 165.535 39.840 168.525 ;
        RECT 37.155 159.820 37.535 160.200 ;
        RECT 40.045 159.840 40.425 161.215 ;
        RECT 40.815 160.660 41.130 171.710 ;
        RECT 41.830 170.405 42.120 172.465 ;
        RECT 44.615 171.005 45.090 174.055 ;
        RECT 49.570 170.915 49.980 174.010 ;
        RECT 48.610 169.255 48.920 169.285 ;
        RECT 41.750 162.550 42.075 164.920 ;
        RECT 43.400 164.595 43.800 168.560 ;
        RECT 42.485 158.810 42.830 161.270 ;
        RECT 44.120 160.490 44.445 163.255 ;
        RECT 45.105 162.525 45.510 165.855 ;
        RECT 48.610 163.155 48.925 169.255 ;
        RECT 49.755 159.550 50.125 168.650 ;
        RECT 50.700 160.615 50.990 172.450 ;
        RECT 54.150 170.890 54.560 173.985 ;
        RECT 58.605 170.345 58.915 172.860 ;
        RECT 51.595 163.110 51.925 169.305 ;
        RECT 54.515 162.580 54.955 165.855 ;
        RECT 56.895 164.595 57.420 168.535 ;
        RECT 56.055 160.490 56.380 163.255 ;
        RECT 58.570 162.585 58.985 164.975 ;
        RECT 59.600 161.145 59.915 171.830 ;
        RECT 60.930 165.535 61.415 168.545 ;
        RECT 62.110 161.160 62.440 171.855 ;
        RECT 60.300 159.755 60.635 161.105 ;
        RECT -78.245 140.890 -77.930 151.940 ;
        RECT -74.410 151.235 -74.010 154.285 ;
        RECT -69.490 151.145 -69.080 154.240 ;
        RECT -64.910 151.120 -64.500 154.215 ;
        RECT -76.575 139.040 -76.230 141.500 ;
        RECT -59.460 141.375 -59.145 152.060 ;
        RECT -55.770 144.170 -55.355 146.985 ;
        RECT -55.030 145.755 -54.645 147.650 ;
        RECT -27.920 140.970 -27.605 152.020 ;
        RECT -24.085 151.315 -23.685 154.365 ;
        RECT -19.165 151.225 -18.755 154.320 ;
        RECT -14.585 151.200 -14.175 154.295 ;
        RECT -26.250 139.120 -25.905 141.580 ;
        RECT -9.135 141.455 -8.820 152.140 ;
        RECT -3.950 144.245 -3.500 148.405 ;
        RECT -2.250 147.225 -1.725 147.665 ;
        RECT 0.015 143.930 0.370 157.720 ;
        RECT 63.360 157.090 63.810 167.355 ;
        RECT 1.640 144.785 2.000 156.120 ;
        RECT 64.525 155.550 65.010 164.435 ;
        RECT 70.830 155.175 71.235 166.705 ;
        RECT 72.905 157.075 73.295 168.175 ;
        RECT 76.675 160.625 77.030 171.710 ;
        RECT 80.420 170.350 80.710 172.410 ;
        RECT 83.190 170.950 83.690 174.000 ;
        RECT 88.160 170.860 88.570 173.955 ;
        RECT 87.200 169.200 87.510 169.230 ;
        RECT 78.000 165.480 78.470 168.470 ;
        RECT 80.350 162.495 80.665 164.865 ;
        RECT 81.970 164.540 82.390 168.505 ;
        RECT 78.635 159.785 79.015 161.160 ;
        RECT 81.075 158.755 81.420 161.215 ;
        RECT 82.710 160.435 83.035 163.200 ;
        RECT 83.695 162.470 84.100 165.800 ;
        RECT 87.200 163.100 87.515 169.200 ;
        RECT 88.345 159.495 88.715 168.595 ;
        RECT 89.290 160.560 89.580 172.395 ;
        RECT 92.740 170.835 93.150 173.930 ;
        RECT 97.195 170.290 97.505 172.805 ;
        RECT 101.445 171.990 101.825 172.370 ;
        RECT 103.575 171.990 103.955 172.370 ;
        RECT 90.185 163.055 90.515 169.250 ;
        RECT 93.090 162.525 93.545 165.800 ;
        RECT 95.450 164.540 95.995 168.480 ;
        RECT 99.505 165.480 99.940 168.490 ;
        RECT 94.645 160.435 94.970 163.200 ;
        RECT 97.160 162.530 97.575 164.920 ;
        RECT 100.700 161.105 101.030 171.800 ;
        RECT 102.135 165.440 102.520 171.225 ;
        RECT 98.890 159.700 99.225 161.050 ;
        RECT 102.495 160.685 102.920 164.960 ;
        RECT 104.195 162.450 104.495 169.490 ;
        RECT 101.155 159.775 101.535 160.155 ;
        RECT 103.350 159.760 103.730 160.140 ;
        RECT 107.220 159.700 107.510 169.480 ;
        RECT 109.070 161.935 109.370 168.745 ;
        RECT 109.860 162.530 110.170 172.570 ;
        RECT 119.050 170.815 119.430 171.195 ;
        RECT 110.655 162.460 110.955 169.290 ;
        RECT 113.230 161.720 113.510 164.755 ;
        RECT 115.980 161.675 116.280 168.830 ;
        RECT 119.655 162.450 119.955 169.490 ;
        RECT 118.950 160.640 119.330 161.020 ;
        RECT 122.680 160.235 122.970 169.480 ;
        RECT 124.530 161.935 124.830 168.745 ;
        RECT 125.320 162.530 125.630 171.265 ;
        RECT 126.115 162.460 126.415 169.290 ;
        RECT 128.690 161.720 128.970 164.755 ;
        RECT 131.440 161.675 131.740 168.830 ;
        RECT 168.335 160.695 168.650 171.745 ;
        RECT 172.170 171.040 172.570 174.090 ;
        RECT 177.090 170.950 177.500 174.045 ;
        RECT 181.670 170.925 182.080 174.020 ;
        RECT 170.005 158.845 170.350 161.305 ;
        RECT 187.120 161.180 187.435 171.865 ;
        RECT 192.305 163.970 192.755 168.130 ;
        RECT 201.700 167.685 202.080 168.065 ;
        RECT 194.005 166.950 194.530 167.390 ;
        RECT 201.690 166.935 202.070 167.315 ;
        RECT 5.290 147.995 5.670 148.375 ;
        RECT 5.280 147.245 5.660 147.625 ;
        RECT 5.325 146.560 5.705 146.940 ;
        RECT 5.290 145.890 5.670 146.270 ;
        RECT 6.005 142.815 6.305 149.855 ;
        RECT 7.125 142.210 7.425 149.140 ;
        RECT 7.780 143.570 8.080 147.630 ;
        RECT 8.435 142.810 8.735 149.160 ;
        RECT 9.030 144.685 9.350 149.845 ;
        RECT 9.750 142.840 10.045 149.665 ;
        RECT 10.880 142.300 11.180 149.110 ;
        RECT 11.670 142.895 11.980 149.085 ;
        RECT 12.465 142.825 12.765 149.655 ;
        RECT 13.590 142.210 13.890 149.150 ;
        RECT 14.270 143.555 14.550 147.645 ;
        RECT 15.040 142.085 15.320 145.120 ;
        RECT 15.800 142.785 16.105 149.145 ;
        RECT 16.650 142.785 16.950 149.605 ;
        RECT 17.790 142.040 18.090 149.195 ;
        RECT 18.455 147.995 18.835 148.375 ;
        RECT 20.725 147.995 21.105 148.400 ;
        RECT 18.460 147.245 18.840 147.625 ;
        RECT 20.730 147.245 21.110 147.650 ;
        RECT 18.460 146.230 18.840 146.610 ;
        RECT 20.245 144.810 20.565 146.940 ;
        RECT 18.675 141.520 19.055 144.540 ;
        RECT 20.855 143.970 21.135 146.375 ;
        RECT 21.465 142.815 21.765 149.855 ;
        RECT 22.585 142.210 22.885 149.140 ;
        RECT 23.240 143.570 23.540 147.630 ;
        RECT 23.895 142.810 24.195 149.160 ;
        RECT 24.490 144.685 24.815 149.845 ;
        RECT 25.210 142.840 25.505 149.665 ;
        RECT 26.340 142.300 26.640 149.110 ;
        RECT 27.130 142.895 27.440 149.085 ;
        RECT 27.925 142.825 28.225 149.655 ;
        RECT 29.050 142.210 29.350 149.150 ;
        RECT 29.730 143.555 30.010 147.645 ;
        RECT 30.500 142.085 30.780 145.120 ;
        RECT 31.260 142.785 31.580 149.145 ;
        RECT 32.110 142.785 32.410 149.605 ;
        RECT 33.250 142.040 33.550 149.195 ;
        RECT 34.190 147.995 34.550 149.825 ;
        RECT 33.885 144.185 34.265 144.565 ;
        RECT 34.590 140.070 34.950 146.630 ;
        RECT 35.730 144.820 36.055 146.685 ;
        RECT 36.370 146.475 36.785 149.825 ;
        RECT 36.395 141.475 36.855 146.160 ;
        RECT 37.180 144.020 37.630 152.840 ;
        RECT 38.040 141.645 38.395 151.950 ;
        RECT 38.705 147.250 39.050 148.305 ;
        RECT 39.365 145.845 39.795 148.835 ;
        RECT 37.110 140.130 37.490 140.510 ;
        RECT 40.000 140.150 40.380 141.525 ;
        RECT 40.770 140.970 41.085 152.020 ;
        RECT 41.785 150.715 42.075 152.775 ;
        RECT 44.570 151.315 45.045 154.365 ;
        RECT 49.525 151.225 49.935 154.320 ;
        RECT 48.565 149.565 48.875 149.595 ;
        RECT 41.705 142.860 42.030 145.230 ;
        RECT 43.355 144.905 43.755 148.870 ;
        RECT 42.440 139.120 42.785 141.580 ;
        RECT 44.075 140.800 44.400 143.565 ;
        RECT 45.060 142.835 45.465 146.165 ;
        RECT 48.565 143.465 48.880 149.565 ;
        RECT 49.710 139.860 50.080 148.960 ;
        RECT 50.655 140.925 50.945 152.760 ;
        RECT 54.105 151.200 54.515 154.295 ;
        RECT 58.560 150.655 58.870 153.170 ;
        RECT 51.550 143.420 51.880 149.615 ;
        RECT 54.470 142.890 54.910 146.165 ;
        RECT 56.850 144.905 57.375 148.845 ;
        RECT 56.010 140.800 56.335 143.565 ;
        RECT 58.525 142.895 58.940 145.285 ;
        RECT 59.555 141.455 59.870 152.140 ;
        RECT 60.885 145.845 61.370 148.855 ;
        RECT 62.065 141.470 62.395 152.165 ;
        RECT 60.255 140.065 60.590 141.415 ;
        RECT -78.185 121.085 -77.870 132.135 ;
        RECT -74.350 131.430 -73.950 134.480 ;
        RECT -69.430 131.340 -69.020 134.435 ;
        RECT -64.850 131.315 -64.440 134.410 ;
        RECT -76.515 119.235 -76.170 121.695 ;
        RECT -59.400 121.570 -59.085 132.255 ;
        RECT -55.710 124.365 -55.295 127.180 ;
        RECT -54.970 125.950 -54.585 127.845 ;
        RECT -27.860 121.165 -27.545 132.215 ;
        RECT -24.025 131.510 -23.625 134.560 ;
        RECT -19.105 131.420 -18.695 134.515 ;
        RECT -14.525 131.395 -14.115 134.490 ;
        RECT -26.190 119.315 -25.845 121.775 ;
        RECT -9.075 121.650 -8.760 132.335 ;
        RECT -3.890 124.440 -3.440 128.600 ;
        RECT -2.190 127.420 -1.665 127.860 ;
        RECT 0.015 124.165 0.370 138.220 ;
        RECT 63.360 137.590 63.810 147.705 ;
        RECT 1.640 124.970 2.000 136.620 ;
        RECT 64.525 136.050 65.010 144.805 ;
        RECT 71.130 135.425 71.535 146.955 ;
        RECT 73.205 137.325 73.595 148.425 ;
        RECT 76.475 140.900 76.830 151.985 ;
        RECT 80.220 150.625 80.510 152.685 ;
        RECT 82.990 151.225 83.490 154.275 ;
        RECT 87.960 151.135 88.370 154.230 ;
        RECT 87.000 149.475 87.310 149.505 ;
        RECT 77.800 145.755 78.270 148.745 ;
        RECT 80.150 142.770 80.465 145.140 ;
        RECT 81.770 144.815 82.190 148.780 ;
        RECT 78.435 140.060 78.815 141.435 ;
        RECT 80.875 139.030 81.220 141.490 ;
        RECT 82.510 140.710 82.835 143.475 ;
        RECT 83.495 142.745 83.900 146.075 ;
        RECT 87.000 143.375 87.315 149.475 ;
        RECT 88.145 139.770 88.515 148.870 ;
        RECT 89.090 140.835 89.380 152.670 ;
        RECT 92.540 151.110 92.950 154.205 ;
        RECT 96.995 150.565 97.305 153.080 ;
        RECT 101.245 152.265 101.625 152.645 ;
        RECT 103.375 152.265 103.755 152.645 ;
        RECT 89.985 143.330 90.315 149.525 ;
        RECT 92.890 142.800 93.345 146.075 ;
        RECT 95.250 144.815 95.795 148.755 ;
        RECT 99.305 145.755 99.740 148.765 ;
        RECT 94.445 140.710 94.770 143.475 ;
        RECT 96.960 142.805 97.375 145.195 ;
        RECT 100.500 141.380 100.830 152.075 ;
        RECT 101.935 145.715 102.320 151.500 ;
        RECT 98.690 139.975 99.025 141.325 ;
        RECT 102.295 140.960 102.720 145.235 ;
        RECT 103.995 142.725 104.295 149.765 ;
        RECT 105.115 142.120 105.415 149.050 ;
        RECT 106.425 142.720 106.725 149.070 ;
        RECT 100.955 140.050 101.335 140.430 ;
        RECT 103.150 140.035 103.530 140.415 ;
        RECT 107.020 139.975 107.310 149.755 ;
        RECT 107.740 142.750 108.035 149.575 ;
        RECT 108.870 142.210 109.170 149.020 ;
        RECT 109.660 142.805 109.970 152.845 ;
        RECT 118.850 151.090 119.230 151.470 ;
        RECT 110.455 142.735 110.755 149.565 ;
        RECT 111.580 142.120 111.880 149.060 ;
        RECT 113.030 141.995 113.310 145.030 ;
        RECT 113.790 142.695 114.070 149.055 ;
        RECT 114.640 142.695 114.940 149.515 ;
        RECT 115.780 141.950 116.080 149.105 ;
        RECT 116.425 146.140 116.805 146.520 ;
        RECT 116.425 144.085 116.805 144.465 ;
        RECT 118.275 143.965 118.590 148.290 ;
        RECT 118.885 146.040 119.165 147.570 ;
        RECT 119.455 142.725 119.755 149.765 ;
        RECT 120.575 142.120 120.875 149.050 ;
        RECT 121.230 143.480 121.530 147.540 ;
        RECT 121.885 142.720 122.185 149.070 ;
        RECT 118.750 140.915 119.130 141.295 ;
        RECT 122.480 140.510 122.770 149.755 ;
        RECT 123.200 142.750 123.495 149.575 ;
        RECT 124.330 142.210 124.630 149.020 ;
        RECT 125.120 142.805 125.430 151.540 ;
        RECT 125.915 142.735 126.215 149.565 ;
        RECT 127.040 142.120 127.340 149.060 ;
        RECT 127.720 143.465 128.000 147.555 ;
        RECT 128.490 141.995 128.770 145.030 ;
        RECT 129.250 142.695 129.530 149.055 ;
        RECT 130.100 142.695 130.400 149.515 ;
        RECT 131.240 141.950 131.540 149.105 ;
        RECT 133.280 147.845 133.655 156.045 ;
        RECT 135.025 147.040 135.325 158.035 ;
        RECT 136.490 145.975 136.870 156.230 ;
        RECT 137.360 143.820 137.795 157.395 ;
        RECT 193.065 156.640 193.580 166.690 ;
        RECT 201.735 166.250 202.115 166.630 ;
        RECT 194.750 155.285 195.335 166.065 ;
        RECT 201.700 165.580 202.080 165.960 ;
        RECT 202.415 162.505 202.715 169.545 ;
        RECT 203.535 161.900 203.835 168.830 ;
        RECT 204.190 163.260 204.490 167.320 ;
        RECT 204.845 162.500 205.145 168.850 ;
        RECT 205.440 164.375 205.760 169.535 ;
        RECT 206.160 162.530 206.455 169.355 ;
        RECT 207.290 161.990 207.590 168.800 ;
        RECT 208.080 162.585 208.390 168.775 ;
        RECT 208.875 162.515 209.175 169.345 ;
        RECT 210.000 161.900 210.300 168.840 ;
        RECT 210.680 163.245 210.960 167.335 ;
        RECT 211.450 161.775 211.730 164.810 ;
        RECT 212.210 162.475 212.515 168.835 ;
        RECT 213.060 162.475 213.360 169.295 ;
        RECT 214.200 161.730 214.500 168.885 ;
        RECT 214.865 167.685 215.245 168.065 ;
        RECT 217.135 167.685 217.515 168.090 ;
        RECT 214.870 166.935 215.250 167.315 ;
        RECT 217.140 166.935 217.520 167.340 ;
        RECT 214.870 165.920 215.250 166.300 ;
        RECT 216.655 164.500 216.975 166.630 ;
        RECT 215.085 161.210 215.465 164.230 ;
        RECT 217.265 163.660 217.545 166.065 ;
        RECT 217.875 162.505 218.175 169.545 ;
        RECT 218.995 161.900 219.295 168.830 ;
        RECT 219.650 163.260 219.950 167.320 ;
        RECT 220.305 162.500 220.605 168.850 ;
        RECT 220.900 164.375 221.225 169.535 ;
        RECT 221.620 162.530 221.915 169.355 ;
        RECT 222.750 161.990 223.050 168.800 ;
        RECT 223.540 162.585 223.850 168.775 ;
        RECT 224.335 162.515 224.635 169.345 ;
        RECT 225.460 161.900 225.760 168.840 ;
        RECT 226.140 163.245 226.420 167.335 ;
        RECT 226.910 161.775 227.190 164.810 ;
        RECT 227.670 162.475 227.990 168.835 ;
        RECT 228.520 162.475 228.820 169.295 ;
        RECT 229.660 161.730 229.960 168.885 ;
        RECT 230.600 167.685 230.960 169.515 ;
        RECT 230.295 163.875 230.675 164.255 ;
        RECT 231.000 159.760 231.360 166.320 ;
        RECT 232.140 164.510 232.465 166.375 ;
        RECT 232.780 166.165 233.195 169.515 ;
        RECT 232.805 161.165 233.265 165.850 ;
        RECT 233.590 163.710 234.040 172.530 ;
        RECT 234.450 161.335 234.805 171.640 ;
        RECT 235.115 166.940 235.460 167.995 ;
        RECT 235.775 165.535 236.205 168.525 ;
        RECT 233.520 159.820 233.900 160.200 ;
        RECT 236.410 159.840 236.790 161.215 ;
        RECT 237.180 160.660 237.495 171.710 ;
        RECT 238.195 170.405 238.485 172.465 ;
        RECT 240.980 171.005 241.455 174.055 ;
        RECT 245.935 170.915 246.345 174.010 ;
        RECT 244.975 169.255 245.285 169.285 ;
        RECT 238.115 162.550 238.440 164.920 ;
        RECT 239.765 164.595 240.165 168.560 ;
        RECT 238.850 158.810 239.195 161.270 ;
        RECT 240.485 160.490 240.810 163.255 ;
        RECT 241.470 162.525 241.875 165.855 ;
        RECT 244.975 163.155 245.290 169.255 ;
        RECT 246.120 159.550 246.490 168.650 ;
        RECT 247.065 160.615 247.355 172.450 ;
        RECT 250.515 170.890 250.925 173.985 ;
        RECT 254.970 170.345 255.280 172.860 ;
        RECT 247.960 163.110 248.290 169.305 ;
        RECT 250.880 162.580 251.320 165.855 ;
        RECT 253.260 164.595 253.785 168.535 ;
        RECT 252.420 160.490 252.745 163.255 ;
        RECT 254.935 162.585 255.350 164.975 ;
        RECT 255.965 161.145 256.280 171.830 ;
        RECT 257.295 165.535 257.780 168.545 ;
        RECT 258.475 161.160 258.805 171.855 ;
        RECT 256.665 159.755 257.000 161.105 ;
        RECT 168.250 140.980 168.565 152.030 ;
        RECT 172.085 151.325 172.485 154.375 ;
        RECT 177.005 151.235 177.415 154.330 ;
        RECT 181.585 151.210 181.995 154.305 ;
        RECT 169.920 139.130 170.265 141.590 ;
        RECT 187.035 141.465 187.350 152.150 ;
        RECT 192.220 144.255 192.670 148.415 ;
        RECT 193.920 147.235 194.445 147.675 ;
        RECT 5.480 128.285 5.860 128.665 ;
        RECT 5.470 127.535 5.850 127.915 ;
        RECT 5.515 126.850 5.895 127.230 ;
        RECT 5.480 126.180 5.860 126.560 ;
        RECT 6.195 123.105 6.495 130.145 ;
        RECT 7.315 122.500 7.615 129.430 ;
        RECT 7.970 123.860 8.270 127.920 ;
        RECT 8.625 123.100 8.925 129.450 ;
        RECT 9.220 124.975 9.540 130.135 ;
        RECT 9.940 123.130 10.235 129.955 ;
        RECT 11.070 122.590 11.370 129.400 ;
        RECT 11.860 123.185 12.170 129.375 ;
        RECT 12.655 123.115 12.955 129.945 ;
        RECT 13.780 122.500 14.080 129.440 ;
        RECT 14.460 123.845 14.740 127.935 ;
        RECT 15.230 122.375 15.510 125.410 ;
        RECT 15.990 123.075 16.295 129.435 ;
        RECT 16.840 123.075 17.140 129.895 ;
        RECT 17.980 122.330 18.280 129.485 ;
        RECT 18.645 128.285 19.025 128.665 ;
        RECT 20.915 128.285 21.295 128.690 ;
        RECT 18.650 127.535 19.030 127.915 ;
        RECT 20.920 127.535 21.300 127.940 ;
        RECT 18.650 126.520 19.030 126.900 ;
        RECT 20.435 125.100 20.755 127.230 ;
        RECT 18.865 121.810 19.245 124.830 ;
        RECT 21.045 124.260 21.325 126.665 ;
        RECT 21.655 123.105 21.955 130.145 ;
        RECT 22.775 122.500 23.075 129.430 ;
        RECT 23.430 123.860 23.730 127.920 ;
        RECT 24.085 123.100 24.385 129.450 ;
        RECT 24.680 124.975 25.005 130.135 ;
        RECT 25.400 123.130 25.695 129.955 ;
        RECT 26.530 122.590 26.830 129.400 ;
        RECT 27.320 123.185 27.630 129.375 ;
        RECT 28.115 123.115 28.415 129.945 ;
        RECT 29.240 122.500 29.540 129.440 ;
        RECT 29.920 123.845 30.200 127.935 ;
        RECT 30.690 122.375 30.970 125.410 ;
        RECT 31.450 123.075 31.770 129.435 ;
        RECT 32.300 123.075 32.600 129.895 ;
        RECT 33.440 122.330 33.740 129.485 ;
        RECT 34.380 128.285 34.740 130.115 ;
        RECT 34.075 124.475 34.455 124.855 ;
        RECT 34.780 120.360 35.140 126.920 ;
        RECT 35.920 125.110 36.245 126.975 ;
        RECT 36.560 126.765 36.975 130.115 ;
        RECT 36.585 121.765 37.045 126.450 ;
        RECT 37.370 124.310 37.820 133.130 ;
        RECT 38.230 121.935 38.585 132.240 ;
        RECT 38.895 127.540 39.240 128.595 ;
        RECT 39.555 126.135 39.985 129.125 ;
        RECT 37.300 120.420 37.680 120.800 ;
        RECT 40.190 120.440 40.570 121.815 ;
        RECT 40.960 121.260 41.275 132.310 ;
        RECT 41.975 131.005 42.265 133.065 ;
        RECT 44.760 131.605 45.235 134.655 ;
        RECT 49.715 131.515 50.125 134.610 ;
        RECT 48.755 129.855 49.065 129.885 ;
        RECT 41.895 123.150 42.220 125.520 ;
        RECT 43.545 125.195 43.945 129.160 ;
        RECT 42.630 119.410 42.975 121.870 ;
        RECT 44.265 121.090 44.590 123.855 ;
        RECT 45.250 123.125 45.655 126.455 ;
        RECT 48.755 123.755 49.070 129.855 ;
        RECT 49.900 120.150 50.270 129.250 ;
        RECT 50.845 121.215 51.135 133.050 ;
        RECT 54.295 131.490 54.705 134.585 ;
        RECT 58.750 130.945 59.060 133.460 ;
        RECT 51.740 123.710 52.070 129.905 ;
        RECT 54.660 123.180 55.100 126.455 ;
        RECT 57.040 125.195 57.565 129.135 ;
        RECT 56.200 121.090 56.525 123.855 ;
        RECT 58.715 123.185 59.130 125.575 ;
        RECT 59.745 121.745 60.060 132.430 ;
        RECT 61.075 126.135 61.560 129.145 ;
        RECT 62.255 121.760 62.585 132.455 ;
        RECT 60.445 120.355 60.780 121.705 ;
        RECT -78.255 101.315 -77.940 112.365 ;
        RECT -74.420 111.660 -74.020 114.710 ;
        RECT -69.500 111.570 -69.090 114.665 ;
        RECT -64.920 111.545 -64.510 114.640 ;
        RECT -76.585 99.465 -76.240 101.925 ;
        RECT -59.470 101.800 -59.155 112.485 ;
        RECT -55.780 104.595 -55.365 107.410 ;
        RECT -55.040 106.180 -54.655 108.075 ;
        RECT -27.930 101.395 -27.615 112.445 ;
        RECT -24.095 111.740 -23.695 114.790 ;
        RECT -19.175 111.650 -18.765 114.745 ;
        RECT -14.595 111.625 -14.185 114.720 ;
        RECT -26.260 99.545 -25.915 102.005 ;
        RECT -9.145 101.880 -8.830 112.565 ;
        RECT -3.960 104.670 -3.510 108.830 ;
        RECT -2.260 107.650 -1.735 108.090 ;
        RECT 0.225 104.390 0.580 118.180 ;
        RECT 63.570 117.550 64.020 128.050 ;
        RECT 1.850 105.245 2.210 116.580 ;
        RECT 64.735 116.010 65.220 125.250 ;
        RECT 71.150 115.765 71.555 127.295 ;
        RECT 73.225 117.665 73.615 128.765 ;
        RECT 76.630 121.255 76.985 132.340 ;
        RECT 80.375 130.980 80.665 133.040 ;
        RECT 83.145 131.580 83.645 134.630 ;
        RECT 88.115 131.490 88.525 134.585 ;
        RECT 87.155 129.830 87.465 129.860 ;
        RECT 77.955 126.110 78.425 129.100 ;
        RECT 80.305 123.125 80.620 125.495 ;
        RECT 81.925 125.170 82.345 129.135 ;
        RECT 78.590 120.415 78.970 121.790 ;
        RECT 81.030 119.385 81.375 121.845 ;
        RECT 82.665 121.065 82.990 123.830 ;
        RECT 83.650 123.100 84.055 126.430 ;
        RECT 87.155 123.730 87.470 129.830 ;
        RECT 88.300 120.125 88.670 129.225 ;
        RECT 89.245 121.190 89.535 133.025 ;
        RECT 92.695 131.465 93.105 134.560 ;
        RECT 97.150 130.920 97.460 133.435 ;
        RECT 101.400 132.620 101.780 133.000 ;
        RECT 103.530 132.620 103.910 133.000 ;
        RECT 90.140 123.685 90.470 129.880 ;
        RECT 93.045 123.155 93.500 126.430 ;
        RECT 95.405 125.170 95.950 129.110 ;
        RECT 99.460 126.110 99.895 129.120 ;
        RECT 94.600 121.065 94.925 123.830 ;
        RECT 97.115 123.160 97.530 125.550 ;
        RECT 100.655 121.735 100.985 132.430 ;
        RECT 102.090 126.070 102.475 131.855 ;
        RECT 98.845 120.330 99.180 121.680 ;
        RECT 102.450 121.315 102.875 125.590 ;
        RECT 104.150 123.080 104.450 130.120 ;
        RECT 105.270 122.475 105.570 129.405 ;
        RECT 106.580 123.075 106.880 129.425 ;
        RECT 101.110 120.405 101.490 120.785 ;
        RECT 103.305 120.390 103.685 120.770 ;
        RECT 107.175 120.330 107.465 130.110 ;
        RECT 107.895 123.105 108.190 129.930 ;
        RECT 109.025 122.565 109.325 129.375 ;
        RECT 109.815 123.160 110.125 133.200 ;
        RECT 119.005 131.445 119.385 131.825 ;
        RECT 110.610 123.090 110.910 129.920 ;
        RECT 111.735 122.475 112.035 129.415 ;
        RECT 113.185 122.350 113.465 125.385 ;
        RECT 113.945 123.050 114.225 129.410 ;
        RECT 114.795 123.050 115.095 129.870 ;
        RECT 115.935 122.305 116.235 129.460 ;
        RECT 116.580 126.495 116.960 126.875 ;
        RECT 116.580 124.440 116.960 124.820 ;
        RECT 118.430 124.320 118.745 128.645 ;
        RECT 119.040 126.395 119.320 127.925 ;
        RECT 119.610 123.080 119.910 130.120 ;
        RECT 120.730 122.475 121.030 129.405 ;
        RECT 121.385 123.835 121.685 127.895 ;
        RECT 122.040 123.075 122.340 129.425 ;
        RECT 118.905 121.270 119.285 121.650 ;
        RECT 122.635 120.865 122.925 130.110 ;
        RECT 123.355 123.105 123.650 129.930 ;
        RECT 124.485 122.565 124.785 129.375 ;
        RECT 125.275 123.160 125.585 131.895 ;
        RECT 126.070 123.090 126.370 129.920 ;
        RECT 127.195 122.475 127.495 129.415 ;
        RECT 127.875 123.820 128.155 127.910 ;
        RECT 128.645 122.350 128.925 125.385 ;
        RECT 129.405 123.050 129.685 129.410 ;
        RECT 130.255 123.050 130.555 129.870 ;
        RECT 131.395 122.305 131.695 129.460 ;
        RECT 133.580 128.095 133.955 136.295 ;
        RECT 135.325 127.290 135.625 138.285 ;
        RECT 136.490 126.330 136.870 136.585 ;
        RECT 137.360 124.175 137.795 137.750 ;
        RECT 193.065 136.950 193.580 147.000 ;
        RECT 194.750 135.595 195.335 146.375 ;
        RECT 196.380 143.930 196.735 157.720 ;
        RECT 259.725 157.090 260.175 167.355 ;
        RECT 198.005 144.785 198.365 156.120 ;
        RECT 260.890 155.550 261.375 164.435 ;
        RECT 267.195 155.175 267.600 166.705 ;
        RECT 269.270 157.075 269.660 168.175 ;
        RECT 273.040 160.625 273.395 171.710 ;
        RECT 276.785 170.350 277.075 172.410 ;
        RECT 279.555 170.950 280.055 174.000 ;
        RECT 284.525 170.860 284.935 173.955 ;
        RECT 283.565 169.200 283.875 169.230 ;
        RECT 274.365 165.480 274.835 168.470 ;
        RECT 276.715 162.495 277.030 164.865 ;
        RECT 278.335 164.540 278.755 168.505 ;
        RECT 275.000 159.785 275.380 161.160 ;
        RECT 277.440 158.755 277.785 161.215 ;
        RECT 279.075 160.435 279.400 163.200 ;
        RECT 280.060 162.470 280.465 165.800 ;
        RECT 283.565 163.100 283.880 169.200 ;
        RECT 284.710 159.495 285.080 168.595 ;
        RECT 285.655 160.560 285.945 172.395 ;
        RECT 289.105 170.835 289.515 173.930 ;
        RECT 293.560 170.290 293.870 172.805 ;
        RECT 297.810 171.990 298.190 172.370 ;
        RECT 299.940 171.990 300.320 172.370 ;
        RECT 286.550 163.055 286.880 169.250 ;
        RECT 289.455 162.525 289.910 165.800 ;
        RECT 291.815 164.540 292.360 168.480 ;
        RECT 295.870 165.480 296.305 168.490 ;
        RECT 291.010 160.435 291.335 163.200 ;
        RECT 293.525 162.530 293.940 164.920 ;
        RECT 297.065 161.105 297.395 171.800 ;
        RECT 298.500 165.440 298.885 171.225 ;
        RECT 295.255 159.700 295.590 161.050 ;
        RECT 298.860 160.685 299.285 164.960 ;
        RECT 300.560 162.450 300.860 169.490 ;
        RECT 301.680 161.845 301.980 168.775 ;
        RECT 302.990 162.445 303.290 168.795 ;
        RECT 297.520 159.775 297.900 160.155 ;
        RECT 299.715 159.760 300.095 160.140 ;
        RECT 303.585 159.700 303.875 169.480 ;
        RECT 304.305 162.475 304.600 169.300 ;
        RECT 305.435 161.935 305.735 168.745 ;
        RECT 306.225 162.530 306.535 172.570 ;
        RECT 315.415 170.815 315.795 171.195 ;
        RECT 307.020 162.460 307.320 169.290 ;
        RECT 308.145 161.845 308.445 168.785 ;
        RECT 309.595 161.720 309.875 164.755 ;
        RECT 310.355 162.420 310.635 168.780 ;
        RECT 311.205 162.420 311.505 169.240 ;
        RECT 312.345 161.675 312.645 168.830 ;
        RECT 312.990 165.865 313.370 166.245 ;
        RECT 312.990 163.810 313.370 164.190 ;
        RECT 314.840 163.690 315.155 168.015 ;
        RECT 315.450 165.765 315.730 167.295 ;
        RECT 316.020 162.450 316.320 169.490 ;
        RECT 317.795 163.205 318.095 167.265 ;
        RECT 315.315 160.640 315.695 161.020 ;
        RECT 319.045 160.235 319.335 169.480 ;
        RECT 320.895 161.935 321.195 168.745 ;
        RECT 321.685 162.530 321.995 171.265 ;
        RECT 322.480 162.460 322.780 169.290 ;
        RECT 324.285 163.190 324.565 167.280 ;
        RECT 325.055 161.720 325.335 164.755 ;
        RECT 327.805 161.675 328.105 168.830 ;
        RECT 364.725 160.655 365.040 171.705 ;
        RECT 368.560 171.000 368.960 174.050 ;
        RECT 373.480 170.910 373.890 174.005 ;
        RECT 378.060 170.885 378.470 173.980 ;
        RECT 366.395 158.805 366.740 161.265 ;
        RECT 383.510 161.140 383.825 171.825 ;
        RECT 388.695 163.930 389.145 168.090 ;
        RECT 398.100 167.635 398.480 168.015 ;
        RECT 390.395 166.910 390.920 167.350 ;
        RECT 398.090 166.885 398.470 167.265 ;
        RECT 201.655 147.995 202.035 148.375 ;
        RECT 201.645 147.245 202.025 147.625 ;
        RECT 201.690 146.560 202.070 146.940 ;
        RECT 201.655 145.890 202.035 146.270 ;
        RECT 202.370 142.815 202.670 149.855 ;
        RECT 203.490 142.210 203.790 149.140 ;
        RECT 204.145 143.570 204.445 147.630 ;
        RECT 204.800 142.810 205.100 149.160 ;
        RECT 205.395 144.685 205.715 149.845 ;
        RECT 206.115 142.840 206.410 149.665 ;
        RECT 207.245 142.300 207.545 149.110 ;
        RECT 208.035 142.895 208.345 149.085 ;
        RECT 208.830 142.825 209.130 149.655 ;
        RECT 209.955 142.210 210.255 149.150 ;
        RECT 210.635 143.555 210.915 147.645 ;
        RECT 211.405 142.085 211.685 145.120 ;
        RECT 212.165 142.785 212.470 149.145 ;
        RECT 213.015 142.785 213.315 149.605 ;
        RECT 214.155 142.040 214.455 149.195 ;
        RECT 214.820 147.995 215.200 148.375 ;
        RECT 217.090 147.995 217.470 148.400 ;
        RECT 214.825 147.245 215.205 147.625 ;
        RECT 217.095 147.245 217.475 147.650 ;
        RECT 214.825 146.230 215.205 146.610 ;
        RECT 216.610 144.810 216.930 146.940 ;
        RECT 215.040 141.520 215.420 144.540 ;
        RECT 217.220 143.970 217.500 146.375 ;
        RECT 217.830 142.815 218.130 149.855 ;
        RECT 218.950 142.210 219.250 149.140 ;
        RECT 219.605 143.570 219.905 147.630 ;
        RECT 220.260 142.810 220.560 149.160 ;
        RECT 220.855 144.685 221.180 149.845 ;
        RECT 221.575 142.840 221.870 149.665 ;
        RECT 222.705 142.300 223.005 149.110 ;
        RECT 223.495 142.895 223.805 149.085 ;
        RECT 224.290 142.825 224.590 149.655 ;
        RECT 225.415 142.210 225.715 149.150 ;
        RECT 226.095 143.555 226.375 147.645 ;
        RECT 226.865 142.085 227.145 145.120 ;
        RECT 227.625 142.785 227.945 149.145 ;
        RECT 228.475 142.785 228.775 149.605 ;
        RECT 229.615 142.040 229.915 149.195 ;
        RECT 230.555 147.995 230.915 149.825 ;
        RECT 230.250 144.185 230.630 144.565 ;
        RECT 230.955 140.070 231.315 146.630 ;
        RECT 232.095 144.820 232.420 146.685 ;
        RECT 232.735 146.475 233.150 149.825 ;
        RECT 232.760 141.475 233.220 146.160 ;
        RECT 233.545 144.020 233.995 152.840 ;
        RECT 234.405 141.645 234.760 151.950 ;
        RECT 235.070 147.250 235.415 148.305 ;
        RECT 235.730 145.845 236.160 148.835 ;
        RECT 233.475 140.130 233.855 140.510 ;
        RECT 236.365 140.150 236.745 141.525 ;
        RECT 237.135 140.970 237.450 152.020 ;
        RECT 238.150 150.715 238.440 152.775 ;
        RECT 240.935 151.315 241.410 154.365 ;
        RECT 245.890 151.225 246.300 154.320 ;
        RECT 244.930 149.565 245.240 149.595 ;
        RECT 238.070 142.860 238.395 145.230 ;
        RECT 239.720 144.905 240.120 148.870 ;
        RECT 238.805 139.120 239.150 141.580 ;
        RECT 240.440 140.800 240.765 143.565 ;
        RECT 241.425 142.835 241.830 146.165 ;
        RECT 244.930 143.465 245.245 149.565 ;
        RECT 246.075 139.860 246.445 148.960 ;
        RECT 247.020 140.925 247.310 152.760 ;
        RECT 250.470 151.200 250.880 154.295 ;
        RECT 254.925 150.655 255.235 153.170 ;
        RECT 247.915 143.420 248.245 149.615 ;
        RECT 250.835 142.890 251.275 146.165 ;
        RECT 253.215 144.905 253.740 148.845 ;
        RECT 252.375 140.800 252.700 143.565 ;
        RECT 254.890 142.895 255.305 145.285 ;
        RECT 255.920 141.455 256.235 152.140 ;
        RECT 257.250 145.845 257.735 148.855 ;
        RECT 258.430 141.470 258.760 152.165 ;
        RECT 256.620 140.065 256.955 141.415 ;
        RECT 168.310 121.175 168.625 132.225 ;
        RECT 172.145 131.520 172.545 134.570 ;
        RECT 177.065 131.430 177.475 134.525 ;
        RECT 181.645 131.405 182.055 134.500 ;
        RECT 169.980 119.325 170.325 121.785 ;
        RECT 187.095 121.660 187.410 132.345 ;
        RECT 192.280 124.450 192.730 128.610 ;
        RECT 193.980 127.430 194.505 127.870 ;
        RECT 5.285 108.445 5.665 108.825 ;
        RECT 5.275 107.695 5.655 108.075 ;
        RECT 5.320 107.010 5.700 107.390 ;
        RECT 5.285 106.340 5.665 106.720 ;
        RECT 6.000 103.265 6.300 110.305 ;
        RECT 7.120 102.660 7.420 109.590 ;
        RECT 7.775 104.020 8.075 108.080 ;
        RECT 8.430 103.260 8.730 109.610 ;
        RECT 9.025 105.135 9.345 110.295 ;
        RECT 9.745 103.290 10.040 110.115 ;
        RECT 10.875 102.750 11.175 109.560 ;
        RECT 11.665 103.345 11.975 109.535 ;
        RECT 12.460 103.275 12.760 110.105 ;
        RECT 13.585 102.660 13.885 109.600 ;
        RECT 14.265 104.005 14.545 108.095 ;
        RECT 15.035 102.535 15.315 105.570 ;
        RECT 15.795 103.235 16.100 109.595 ;
        RECT 16.645 103.235 16.945 110.055 ;
        RECT 17.785 102.490 18.085 109.645 ;
        RECT 18.450 108.445 18.830 108.825 ;
        RECT 20.720 108.445 21.100 108.850 ;
        RECT 18.455 107.695 18.835 108.075 ;
        RECT 20.725 107.695 21.105 108.100 ;
        RECT 18.455 106.680 18.835 107.060 ;
        RECT 20.240 105.260 20.560 107.390 ;
        RECT 18.670 101.970 19.050 104.990 ;
        RECT 20.850 104.420 21.130 106.825 ;
        RECT 21.460 103.265 21.760 110.305 ;
        RECT 22.580 102.660 22.880 109.590 ;
        RECT 23.235 104.020 23.535 108.080 ;
        RECT 23.890 103.260 24.190 109.610 ;
        RECT 24.485 105.135 24.810 110.295 ;
        RECT 25.205 103.290 25.500 110.115 ;
        RECT 26.335 102.750 26.635 109.560 ;
        RECT 27.125 103.345 27.435 109.535 ;
        RECT 27.920 103.275 28.220 110.105 ;
        RECT 29.045 102.660 29.345 109.600 ;
        RECT 29.725 104.005 30.005 108.095 ;
        RECT 30.495 102.535 30.775 105.570 ;
        RECT 31.255 103.235 31.575 109.595 ;
        RECT 32.105 103.235 32.405 110.055 ;
        RECT 33.245 102.490 33.545 109.645 ;
        RECT 34.185 108.445 34.545 110.275 ;
        RECT 33.880 104.635 34.260 105.015 ;
        RECT 34.585 100.520 34.945 107.080 ;
        RECT 35.725 105.270 36.050 107.135 ;
        RECT 36.365 106.925 36.780 110.275 ;
        RECT 36.390 101.925 36.850 106.610 ;
        RECT 37.175 104.470 37.625 113.290 ;
        RECT 38.035 102.095 38.390 112.400 ;
        RECT 38.700 107.700 39.045 108.755 ;
        RECT 39.360 106.295 39.790 109.285 ;
        RECT 37.105 100.580 37.485 100.960 ;
        RECT 39.995 100.600 40.375 101.975 ;
        RECT 40.765 101.420 41.080 112.470 ;
        RECT 41.780 111.165 42.070 113.225 ;
        RECT 44.565 111.765 45.040 114.815 ;
        RECT 49.520 111.675 49.930 114.770 ;
        RECT 48.560 110.015 48.870 110.045 ;
        RECT 41.700 103.310 42.025 105.680 ;
        RECT 43.350 105.355 43.750 109.320 ;
        RECT 42.435 99.570 42.780 102.030 ;
        RECT 44.070 101.250 44.395 104.015 ;
        RECT 45.055 103.285 45.460 106.615 ;
        RECT 48.560 103.915 48.875 110.015 ;
        RECT 49.705 100.310 50.075 109.410 ;
        RECT 50.650 101.375 50.940 113.210 ;
        RECT 54.100 111.650 54.510 114.745 ;
        RECT 58.555 111.105 58.865 113.620 ;
        RECT 51.545 103.870 51.875 110.065 ;
        RECT 54.465 103.340 54.905 106.615 ;
        RECT 56.845 105.355 57.370 109.295 ;
        RECT 56.005 101.250 56.330 104.015 ;
        RECT 58.520 103.345 58.935 105.735 ;
        RECT 59.550 101.905 59.865 112.590 ;
        RECT 60.880 106.295 61.365 109.305 ;
        RECT 62.060 101.920 62.390 112.615 ;
        RECT 60.250 100.515 60.585 101.865 ;
        RECT -78.225 81.590 -77.910 92.640 ;
        RECT -74.390 91.935 -73.990 94.985 ;
        RECT -69.470 91.845 -69.060 94.940 ;
        RECT -64.890 91.820 -64.480 94.915 ;
        RECT -76.555 79.740 -76.210 82.200 ;
        RECT -59.440 82.075 -59.125 92.760 ;
        RECT -55.750 84.870 -55.335 87.685 ;
        RECT -55.010 86.455 -54.625 88.350 ;
        RECT -27.900 81.670 -27.585 92.720 ;
        RECT -24.065 92.015 -23.665 95.065 ;
        RECT -19.145 91.925 -18.735 95.020 ;
        RECT -14.565 91.900 -14.155 94.995 ;
        RECT -26.230 79.820 -25.885 82.280 ;
        RECT -9.115 82.155 -8.800 92.840 ;
        RECT -3.930 84.945 -3.480 89.105 ;
        RECT -2.230 87.925 -1.705 88.365 ;
        RECT 0.180 84.600 0.535 98.390 ;
        RECT 63.525 97.760 63.975 108.250 ;
        RECT 1.805 85.505 2.165 96.790 ;
        RECT 64.690 96.220 65.175 105.380 ;
        RECT 71.150 96.030 71.555 107.560 ;
        RECT 73.225 97.930 73.615 109.030 ;
        RECT 76.630 101.460 76.985 112.545 ;
        RECT 80.375 111.185 80.665 113.245 ;
        RECT 83.145 111.785 83.645 114.835 ;
        RECT 88.115 111.695 88.525 114.790 ;
        RECT 87.155 110.035 87.465 110.065 ;
        RECT 77.955 106.315 78.425 109.305 ;
        RECT 80.305 103.330 80.620 105.700 ;
        RECT 81.925 105.375 82.345 109.340 ;
        RECT 78.590 100.620 78.970 101.995 ;
        RECT 81.030 99.590 81.375 102.050 ;
        RECT 82.665 101.270 82.990 104.035 ;
        RECT 83.650 103.305 84.055 106.635 ;
        RECT 87.155 103.935 87.470 110.035 ;
        RECT 88.300 100.330 88.670 109.430 ;
        RECT 89.245 101.395 89.535 113.230 ;
        RECT 92.695 111.670 93.105 114.765 ;
        RECT 97.150 111.125 97.460 113.640 ;
        RECT 101.400 112.825 101.780 113.205 ;
        RECT 103.530 112.825 103.910 113.205 ;
        RECT 90.140 103.890 90.470 110.085 ;
        RECT 93.045 103.360 93.500 106.635 ;
        RECT 95.405 105.375 95.950 109.315 ;
        RECT 99.460 106.315 99.895 109.325 ;
        RECT 94.600 101.270 94.925 104.035 ;
        RECT 97.115 103.365 97.530 105.755 ;
        RECT 100.655 101.940 100.985 112.635 ;
        RECT 102.090 106.275 102.475 112.060 ;
        RECT 98.845 100.535 99.180 101.885 ;
        RECT 102.450 101.520 102.875 105.795 ;
        RECT 104.150 103.285 104.450 110.325 ;
        RECT 105.270 102.680 105.570 109.610 ;
        RECT 106.580 103.280 106.880 109.630 ;
        RECT 101.110 100.610 101.490 100.990 ;
        RECT 103.305 100.595 103.685 100.975 ;
        RECT 107.175 100.535 107.465 110.315 ;
        RECT 107.895 103.310 108.190 110.135 ;
        RECT 109.025 102.770 109.325 109.580 ;
        RECT 109.815 103.365 110.125 113.405 ;
        RECT 119.005 111.650 119.385 112.030 ;
        RECT 110.610 103.295 110.910 110.125 ;
        RECT 111.735 102.680 112.035 109.620 ;
        RECT 113.185 102.555 113.465 105.590 ;
        RECT 113.945 103.255 114.225 109.615 ;
        RECT 114.795 103.255 115.095 110.075 ;
        RECT 115.935 102.510 116.235 109.665 ;
        RECT 116.580 106.700 116.960 107.080 ;
        RECT 116.580 104.645 116.960 105.025 ;
        RECT 118.430 104.525 118.745 108.850 ;
        RECT 119.040 106.600 119.320 108.130 ;
        RECT 119.610 103.285 119.910 110.325 ;
        RECT 120.730 102.680 121.030 109.610 ;
        RECT 121.385 104.040 121.685 108.100 ;
        RECT 122.040 103.280 122.340 109.630 ;
        RECT 118.905 101.475 119.285 101.855 ;
        RECT 122.635 101.070 122.925 110.315 ;
        RECT 123.355 103.310 123.650 110.135 ;
        RECT 124.485 102.770 124.785 109.580 ;
        RECT 125.275 103.365 125.585 112.100 ;
        RECT 126.070 103.295 126.370 110.125 ;
        RECT 127.195 102.680 127.495 109.620 ;
        RECT 127.875 104.025 128.155 108.115 ;
        RECT 128.645 102.555 128.925 105.590 ;
        RECT 129.405 103.255 129.685 109.615 ;
        RECT 130.255 103.255 130.555 110.075 ;
        RECT 131.395 102.510 131.695 109.665 ;
        RECT 133.600 108.435 133.975 116.635 ;
        RECT 135.345 107.630 135.645 118.625 ;
        RECT 136.490 106.535 136.870 116.790 ;
        RECT 137.360 104.380 137.795 117.955 ;
        RECT 193.215 117.235 193.730 127.285 ;
        RECT 194.900 115.880 195.485 126.660 ;
        RECT 196.380 124.165 196.735 138.220 ;
        RECT 259.725 137.590 260.175 147.705 ;
        RECT 198.005 124.970 198.365 136.620 ;
        RECT 260.890 136.050 261.375 144.805 ;
        RECT 267.495 135.425 267.900 146.955 ;
        RECT 269.570 137.325 269.960 148.425 ;
        RECT 272.840 140.900 273.195 151.985 ;
        RECT 276.585 150.625 276.875 152.685 ;
        RECT 279.355 151.225 279.855 154.275 ;
        RECT 284.325 151.135 284.735 154.230 ;
        RECT 283.365 149.475 283.675 149.505 ;
        RECT 274.165 145.755 274.635 148.745 ;
        RECT 276.515 142.770 276.830 145.140 ;
        RECT 278.135 144.815 278.555 148.780 ;
        RECT 274.800 140.060 275.180 141.435 ;
        RECT 277.240 139.030 277.585 141.490 ;
        RECT 278.875 140.710 279.200 143.475 ;
        RECT 279.860 142.745 280.265 146.075 ;
        RECT 283.365 143.375 283.680 149.475 ;
        RECT 284.510 139.770 284.880 148.870 ;
        RECT 285.455 140.835 285.745 152.670 ;
        RECT 288.905 151.110 289.315 154.205 ;
        RECT 293.360 150.565 293.670 153.080 ;
        RECT 297.610 152.265 297.990 152.645 ;
        RECT 299.740 152.265 300.120 152.645 ;
        RECT 286.350 143.330 286.680 149.525 ;
        RECT 289.255 142.800 289.710 146.075 ;
        RECT 291.615 144.815 292.160 148.755 ;
        RECT 295.670 145.755 296.105 148.765 ;
        RECT 290.810 140.710 291.135 143.475 ;
        RECT 293.325 142.805 293.740 145.195 ;
        RECT 296.865 141.380 297.195 152.075 ;
        RECT 298.300 145.715 298.685 151.500 ;
        RECT 295.055 139.975 295.390 141.325 ;
        RECT 298.660 140.960 299.085 145.235 ;
        RECT 300.360 142.725 300.660 149.765 ;
        RECT 301.480 142.120 301.780 149.050 ;
        RECT 302.790 142.720 303.090 149.070 ;
        RECT 297.320 140.050 297.700 140.430 ;
        RECT 299.515 140.035 299.895 140.415 ;
        RECT 303.385 139.975 303.675 149.755 ;
        RECT 304.105 142.750 304.400 149.575 ;
        RECT 305.235 142.210 305.535 149.020 ;
        RECT 306.025 142.805 306.335 152.845 ;
        RECT 315.215 151.090 315.595 151.470 ;
        RECT 306.820 142.735 307.120 149.565 ;
        RECT 307.945 142.120 308.245 149.060 ;
        RECT 309.395 141.995 309.675 145.030 ;
        RECT 310.155 142.695 310.435 149.055 ;
        RECT 311.005 142.695 311.305 149.515 ;
        RECT 312.145 141.950 312.445 149.105 ;
        RECT 312.790 146.140 313.170 146.520 ;
        RECT 312.790 144.085 313.170 144.465 ;
        RECT 314.640 143.965 314.955 148.290 ;
        RECT 315.250 146.040 315.530 147.570 ;
        RECT 315.820 142.725 316.120 149.765 ;
        RECT 316.940 142.120 317.240 149.050 ;
        RECT 317.595 143.480 317.895 147.540 ;
        RECT 318.250 142.720 318.550 149.070 ;
        RECT 315.115 140.915 315.495 141.295 ;
        RECT 318.845 140.510 319.135 149.755 ;
        RECT 319.565 142.750 319.860 149.575 ;
        RECT 320.695 142.210 320.995 149.020 ;
        RECT 321.485 142.805 321.795 151.540 ;
        RECT 322.280 142.735 322.580 149.565 ;
        RECT 323.405 142.120 323.705 149.060 ;
        RECT 324.085 143.465 324.365 147.555 ;
        RECT 324.855 141.995 325.135 145.030 ;
        RECT 325.615 142.695 325.895 149.055 ;
        RECT 326.465 142.695 326.765 149.515 ;
        RECT 327.605 141.950 327.905 149.105 ;
        RECT 329.645 147.845 330.020 156.045 ;
        RECT 331.390 147.040 331.690 158.035 ;
        RECT 332.880 145.935 333.260 156.190 ;
        RECT 333.750 143.780 334.185 157.355 ;
        RECT 389.455 156.600 389.970 166.650 ;
        RECT 398.135 166.200 398.515 166.580 ;
        RECT 391.140 155.245 391.725 166.025 ;
        RECT 398.100 165.530 398.480 165.910 ;
        RECT 398.815 162.455 399.115 169.495 ;
        RECT 399.935 161.850 400.235 168.780 ;
        RECT 400.590 163.210 400.890 167.270 ;
        RECT 401.245 162.450 401.545 168.800 ;
        RECT 401.840 164.325 402.160 169.485 ;
        RECT 402.560 162.480 402.855 169.305 ;
        RECT 403.690 161.940 403.990 168.750 ;
        RECT 404.480 162.535 404.790 168.725 ;
        RECT 405.275 162.465 405.575 169.295 ;
        RECT 406.400 161.850 406.700 168.790 ;
        RECT 407.080 163.195 407.360 167.285 ;
        RECT 407.850 161.725 408.130 164.760 ;
        RECT 408.610 162.425 408.915 168.785 ;
        RECT 409.460 162.425 409.760 169.245 ;
        RECT 410.600 161.680 410.900 168.835 ;
        RECT 411.265 167.635 411.645 168.015 ;
        RECT 413.535 167.635 413.915 168.040 ;
        RECT 411.270 166.885 411.650 167.265 ;
        RECT 413.540 166.885 413.920 167.290 ;
        RECT 411.270 165.870 411.650 166.250 ;
        RECT 413.055 164.450 413.375 166.580 ;
        RECT 411.485 161.160 411.865 164.180 ;
        RECT 413.665 163.610 413.945 166.015 ;
        RECT 414.275 162.455 414.575 169.495 ;
        RECT 415.395 161.850 415.695 168.780 ;
        RECT 416.050 163.210 416.350 167.270 ;
        RECT 416.705 162.450 417.005 168.800 ;
        RECT 417.300 164.325 417.625 169.485 ;
        RECT 418.020 162.480 418.315 169.305 ;
        RECT 419.150 161.940 419.450 168.750 ;
        RECT 419.940 162.535 420.250 168.725 ;
        RECT 420.735 162.465 421.035 169.295 ;
        RECT 421.860 161.850 422.160 168.790 ;
        RECT 422.540 163.195 422.820 167.285 ;
        RECT 423.310 161.725 423.590 164.760 ;
        RECT 424.070 162.425 424.390 168.785 ;
        RECT 424.920 162.425 425.220 169.245 ;
        RECT 426.060 161.680 426.360 168.835 ;
        RECT 427.000 167.635 427.360 169.465 ;
        RECT 426.695 163.825 427.075 164.205 ;
        RECT 427.400 159.710 427.760 166.270 ;
        RECT 428.540 164.460 428.865 166.325 ;
        RECT 429.180 166.115 429.595 169.465 ;
        RECT 429.205 161.115 429.665 165.800 ;
        RECT 429.990 163.660 430.440 172.480 ;
        RECT 430.850 161.285 431.205 171.590 ;
        RECT 431.515 166.890 431.860 167.945 ;
        RECT 432.175 165.485 432.605 168.475 ;
        RECT 429.920 159.770 430.300 160.150 ;
        RECT 432.810 159.790 433.190 161.165 ;
        RECT 433.580 160.610 433.895 171.660 ;
        RECT 434.595 170.355 434.885 172.415 ;
        RECT 437.380 170.955 437.855 174.005 ;
        RECT 442.335 170.865 442.745 173.960 ;
        RECT 441.375 169.205 441.685 169.235 ;
        RECT 434.515 162.500 434.840 164.870 ;
        RECT 436.165 164.545 436.565 168.510 ;
        RECT 435.250 158.760 435.595 161.220 ;
        RECT 436.885 160.440 437.210 163.205 ;
        RECT 437.870 162.475 438.275 165.805 ;
        RECT 441.375 163.105 441.690 169.205 ;
        RECT 442.520 159.500 442.890 168.600 ;
        RECT 443.465 160.565 443.755 172.400 ;
        RECT 446.915 170.840 447.325 173.935 ;
        RECT 451.370 170.295 451.680 172.810 ;
        RECT 444.360 163.060 444.690 169.255 ;
        RECT 447.280 162.530 447.720 165.805 ;
        RECT 449.660 164.545 450.185 168.485 ;
        RECT 448.820 160.440 449.145 163.205 ;
        RECT 451.335 162.535 451.750 164.925 ;
        RECT 452.365 161.095 452.680 171.780 ;
        RECT 453.695 165.485 454.180 168.495 ;
        RECT 454.875 161.110 455.205 171.805 ;
        RECT 453.065 159.705 453.400 161.055 ;
        RECT 364.640 140.940 364.955 151.990 ;
        RECT 368.475 151.285 368.875 154.335 ;
        RECT 373.395 151.195 373.805 154.290 ;
        RECT 377.975 151.170 378.385 154.265 ;
        RECT 366.310 139.090 366.655 141.550 ;
        RECT 383.425 141.425 383.740 152.110 ;
        RECT 388.610 144.215 389.060 148.375 ;
        RECT 390.310 147.195 390.835 147.635 ;
        RECT 201.845 128.285 202.225 128.665 ;
        RECT 201.835 127.535 202.215 127.915 ;
        RECT 201.880 126.850 202.260 127.230 ;
        RECT 201.845 126.180 202.225 126.560 ;
        RECT 202.560 123.105 202.860 130.145 ;
        RECT 203.680 122.500 203.980 129.430 ;
        RECT 204.335 123.860 204.635 127.920 ;
        RECT 204.990 123.100 205.290 129.450 ;
        RECT 205.585 124.975 205.905 130.135 ;
        RECT 206.305 123.130 206.600 129.955 ;
        RECT 207.435 122.590 207.735 129.400 ;
        RECT 208.225 123.185 208.535 129.375 ;
        RECT 209.020 123.115 209.320 129.945 ;
        RECT 210.145 122.500 210.445 129.440 ;
        RECT 210.825 123.845 211.105 127.935 ;
        RECT 211.595 122.375 211.875 125.410 ;
        RECT 212.355 123.075 212.660 129.435 ;
        RECT 213.205 123.075 213.505 129.895 ;
        RECT 214.345 122.330 214.645 129.485 ;
        RECT 215.010 128.285 215.390 128.665 ;
        RECT 217.280 128.285 217.660 128.690 ;
        RECT 215.015 127.535 215.395 127.915 ;
        RECT 217.285 127.535 217.665 127.940 ;
        RECT 215.015 126.520 215.395 126.900 ;
        RECT 216.800 125.100 217.120 127.230 ;
        RECT 215.230 121.810 215.610 124.830 ;
        RECT 217.410 124.260 217.690 126.665 ;
        RECT 218.020 123.105 218.320 130.145 ;
        RECT 219.140 122.500 219.440 129.430 ;
        RECT 219.795 123.860 220.095 127.920 ;
        RECT 220.450 123.100 220.750 129.450 ;
        RECT 221.045 124.975 221.370 130.135 ;
        RECT 221.765 123.130 222.060 129.955 ;
        RECT 222.895 122.590 223.195 129.400 ;
        RECT 223.685 123.185 223.995 129.375 ;
        RECT 224.480 123.115 224.780 129.945 ;
        RECT 225.605 122.500 225.905 129.440 ;
        RECT 226.285 123.845 226.565 127.935 ;
        RECT 227.055 122.375 227.335 125.410 ;
        RECT 227.815 123.075 228.135 129.435 ;
        RECT 228.665 123.075 228.965 129.895 ;
        RECT 229.805 122.330 230.105 129.485 ;
        RECT 230.745 128.285 231.105 130.115 ;
        RECT 230.440 124.475 230.820 124.855 ;
        RECT 231.145 120.360 231.505 126.920 ;
        RECT 232.285 125.110 232.610 126.975 ;
        RECT 232.925 126.765 233.340 130.115 ;
        RECT 232.950 121.765 233.410 126.450 ;
        RECT 233.735 124.310 234.185 133.130 ;
        RECT 234.595 121.935 234.950 132.240 ;
        RECT 235.260 127.540 235.605 128.595 ;
        RECT 235.920 126.135 236.350 129.125 ;
        RECT 233.665 120.420 234.045 120.800 ;
        RECT 236.555 120.440 236.935 121.815 ;
        RECT 237.325 121.260 237.640 132.310 ;
        RECT 238.340 131.005 238.630 133.065 ;
        RECT 241.125 131.605 241.600 134.655 ;
        RECT 246.080 131.515 246.490 134.610 ;
        RECT 245.120 129.855 245.430 129.885 ;
        RECT 238.260 123.150 238.585 125.520 ;
        RECT 239.910 125.195 240.310 129.160 ;
        RECT 238.995 119.410 239.340 121.870 ;
        RECT 240.630 121.090 240.955 123.855 ;
        RECT 241.615 123.125 242.020 126.455 ;
        RECT 245.120 123.755 245.435 129.855 ;
        RECT 246.265 120.150 246.635 129.250 ;
        RECT 247.210 121.215 247.500 133.050 ;
        RECT 250.660 131.490 251.070 134.585 ;
        RECT 255.115 130.945 255.425 133.460 ;
        RECT 248.105 123.710 248.435 129.905 ;
        RECT 251.025 123.180 251.465 126.455 ;
        RECT 253.405 125.195 253.930 129.135 ;
        RECT 252.565 121.090 252.890 123.855 ;
        RECT 255.080 123.185 255.495 125.575 ;
        RECT 256.110 121.745 256.425 132.430 ;
        RECT 257.440 126.135 257.925 129.145 ;
        RECT 258.620 121.760 258.950 132.455 ;
        RECT 256.810 120.355 257.145 121.705 ;
        RECT 168.240 101.405 168.555 112.455 ;
        RECT 172.075 111.750 172.475 114.800 ;
        RECT 176.995 111.660 177.405 114.755 ;
        RECT 181.575 111.635 181.985 114.730 ;
        RECT 169.910 99.555 170.255 102.015 ;
        RECT 187.025 101.890 187.340 112.575 ;
        RECT 192.210 104.680 192.660 108.840 ;
        RECT 193.910 107.660 194.435 108.100 ;
        RECT 5.155 88.735 5.535 89.115 ;
        RECT 5.145 87.985 5.525 88.365 ;
        RECT 5.190 87.300 5.570 87.680 ;
        RECT 5.155 86.630 5.535 87.010 ;
        RECT 5.870 83.555 6.170 90.595 ;
        RECT 6.990 82.950 7.290 89.880 ;
        RECT 7.645 84.310 7.945 88.370 ;
        RECT 8.300 83.550 8.600 89.900 ;
        RECT 8.895 85.425 9.215 90.585 ;
        RECT 9.615 83.580 9.910 90.405 ;
        RECT 10.745 83.040 11.045 89.850 ;
        RECT 11.535 83.635 11.845 89.825 ;
        RECT 12.330 83.565 12.630 90.395 ;
        RECT 13.455 82.950 13.755 89.890 ;
        RECT 14.135 84.295 14.415 88.385 ;
        RECT 14.905 82.825 15.185 85.860 ;
        RECT 15.665 83.525 15.970 89.885 ;
        RECT 16.515 83.525 16.815 90.345 ;
        RECT 17.655 82.780 17.955 89.935 ;
        RECT 18.320 88.735 18.700 89.115 ;
        RECT 20.590 88.735 20.970 89.140 ;
        RECT 18.325 87.985 18.705 88.365 ;
        RECT 20.595 87.985 20.975 88.390 ;
        RECT 18.325 86.970 18.705 87.350 ;
        RECT 20.110 85.550 20.430 87.680 ;
        RECT 18.540 82.260 18.920 85.280 ;
        RECT 20.720 84.710 21.000 87.115 ;
        RECT 21.330 83.555 21.630 90.595 ;
        RECT 22.450 82.950 22.750 89.880 ;
        RECT 23.105 84.310 23.405 88.370 ;
        RECT 23.760 83.550 24.060 89.900 ;
        RECT 24.355 85.425 24.680 90.585 ;
        RECT 25.075 83.580 25.370 90.405 ;
        RECT 26.205 83.040 26.505 89.850 ;
        RECT 26.995 83.635 27.305 89.825 ;
        RECT 27.790 83.565 28.090 90.395 ;
        RECT 28.915 82.950 29.215 89.890 ;
        RECT 29.595 84.295 29.875 88.385 ;
        RECT 30.365 82.825 30.645 85.860 ;
        RECT 31.125 83.525 31.445 89.885 ;
        RECT 31.975 83.525 32.275 90.345 ;
        RECT 33.115 82.780 33.415 89.935 ;
        RECT 34.055 88.735 34.415 90.565 ;
        RECT 33.750 84.925 34.130 85.305 ;
        RECT 34.455 80.810 34.815 87.370 ;
        RECT 35.595 85.560 35.920 87.425 ;
        RECT 36.235 87.215 36.650 90.565 ;
        RECT 36.260 82.215 36.720 86.900 ;
        RECT 37.045 84.760 37.495 93.580 ;
        RECT 37.905 82.385 38.260 92.690 ;
        RECT 38.570 87.990 38.915 89.045 ;
        RECT 39.230 86.585 39.660 89.575 ;
        RECT 36.975 80.870 37.355 81.250 ;
        RECT 39.865 80.890 40.245 82.265 ;
        RECT 40.635 81.710 40.950 92.760 ;
        RECT 41.650 91.455 41.940 93.515 ;
        RECT 44.435 92.055 44.910 95.105 ;
        RECT 49.390 91.965 49.800 95.060 ;
        RECT 48.430 90.305 48.740 90.335 ;
        RECT 41.570 83.600 41.895 85.970 ;
        RECT 43.220 85.645 43.620 89.610 ;
        RECT 42.305 79.860 42.650 82.320 ;
        RECT 43.940 81.540 44.265 84.305 ;
        RECT 44.925 83.575 45.330 86.905 ;
        RECT 48.430 84.205 48.745 90.305 ;
        RECT 49.575 80.600 49.945 89.700 ;
        RECT 50.520 81.665 50.810 93.500 ;
        RECT 53.970 91.940 54.380 95.035 ;
        RECT 58.425 91.395 58.735 93.910 ;
        RECT 51.415 84.160 51.745 90.355 ;
        RECT 54.335 83.630 54.775 86.905 ;
        RECT 56.715 85.645 57.240 89.585 ;
        RECT 55.875 81.540 56.200 84.305 ;
        RECT 58.390 83.635 58.805 86.025 ;
        RECT 59.420 82.195 59.735 92.880 ;
        RECT 60.750 86.585 61.235 89.595 ;
        RECT 61.930 82.210 62.260 92.905 ;
        RECT 60.120 80.805 60.455 82.155 ;
        RECT -78.295 61.760 -77.980 72.810 ;
        RECT -74.460 72.105 -74.060 75.155 ;
        RECT -69.540 72.015 -69.130 75.110 ;
        RECT -64.960 71.990 -64.550 75.085 ;
        RECT -76.625 59.910 -76.280 62.370 ;
        RECT -59.510 62.245 -59.195 72.930 ;
        RECT -55.820 65.040 -55.405 67.855 ;
        RECT -55.080 66.625 -54.695 68.520 ;
        RECT -27.970 61.840 -27.655 72.890 ;
        RECT -24.135 72.185 -23.735 75.235 ;
        RECT -19.215 72.095 -18.805 75.190 ;
        RECT -14.635 72.070 -14.225 75.165 ;
        RECT -26.300 59.990 -25.955 62.450 ;
        RECT -9.185 62.325 -8.870 73.010 ;
        RECT -4.000 65.115 -3.550 69.275 ;
        RECT -2.300 68.095 -1.775 68.535 ;
        RECT -0.125 64.840 0.230 78.760 ;
        RECT 63.220 78.130 63.670 88.395 ;
        RECT 1.500 65.745 1.860 77.160 ;
        RECT 64.385 76.590 64.870 85.475 ;
        RECT 71.050 76.325 71.455 87.855 ;
        RECT 73.125 78.225 73.515 89.325 ;
        RECT 76.550 81.705 76.905 92.790 ;
        RECT 80.295 91.430 80.585 93.490 ;
        RECT 83.065 92.030 83.565 95.080 ;
        RECT 88.035 91.940 88.445 95.035 ;
        RECT 87.075 90.280 87.385 90.310 ;
        RECT 77.875 86.560 78.345 89.550 ;
        RECT 80.225 83.575 80.540 85.945 ;
        RECT 81.845 85.620 82.265 89.585 ;
        RECT 78.510 80.865 78.890 82.240 ;
        RECT 80.950 79.835 81.295 82.295 ;
        RECT 82.585 81.515 82.910 84.280 ;
        RECT 83.570 83.550 83.975 86.880 ;
        RECT 87.075 84.180 87.390 90.280 ;
        RECT 88.220 80.575 88.590 89.675 ;
        RECT 89.165 81.640 89.455 93.475 ;
        RECT 92.615 91.915 93.025 95.010 ;
        RECT 97.070 91.370 97.380 93.885 ;
        RECT 101.320 93.070 101.700 93.450 ;
        RECT 103.450 93.070 103.830 93.450 ;
        RECT 90.060 84.135 90.390 90.330 ;
        RECT 92.965 83.605 93.420 86.880 ;
        RECT 95.325 85.620 95.870 89.560 ;
        RECT 99.380 86.560 99.815 89.570 ;
        RECT 94.520 81.515 94.845 84.280 ;
        RECT 97.035 83.610 97.450 86.000 ;
        RECT 100.575 82.185 100.905 92.880 ;
        RECT 102.010 86.520 102.395 92.305 ;
        RECT 98.765 80.780 99.100 82.130 ;
        RECT 102.370 81.765 102.795 86.040 ;
        RECT 104.070 83.530 104.370 90.570 ;
        RECT 105.190 82.925 105.490 89.855 ;
        RECT 106.500 83.525 106.800 89.875 ;
        RECT 101.030 80.855 101.410 81.235 ;
        RECT 103.225 80.840 103.605 81.220 ;
        RECT 107.095 80.780 107.385 90.560 ;
        RECT 107.815 83.555 108.110 90.380 ;
        RECT 108.945 83.015 109.245 89.825 ;
        RECT 109.735 83.610 110.045 93.650 ;
        RECT 118.925 91.895 119.305 92.275 ;
        RECT 110.530 83.540 110.830 90.370 ;
        RECT 111.655 82.925 111.955 89.865 ;
        RECT 113.105 82.800 113.385 85.835 ;
        RECT 113.865 83.500 114.145 89.860 ;
        RECT 114.715 83.500 115.015 90.320 ;
        RECT 115.855 82.755 116.155 89.910 ;
        RECT 116.500 86.945 116.880 87.325 ;
        RECT 116.500 84.890 116.880 85.270 ;
        RECT 118.350 84.770 118.665 89.095 ;
        RECT 118.960 86.845 119.240 88.375 ;
        RECT 119.530 83.530 119.830 90.570 ;
        RECT 120.650 82.925 120.950 89.855 ;
        RECT 121.305 84.285 121.605 88.345 ;
        RECT 121.960 83.525 122.260 89.875 ;
        RECT 118.825 81.720 119.205 82.100 ;
        RECT 122.555 81.315 122.845 90.560 ;
        RECT 123.275 83.555 123.570 90.380 ;
        RECT 124.405 83.015 124.705 89.825 ;
        RECT 125.195 83.610 125.505 92.345 ;
        RECT 125.990 83.540 126.290 90.370 ;
        RECT 127.115 82.925 127.415 89.865 ;
        RECT 127.795 84.270 128.075 88.360 ;
        RECT 128.565 82.800 128.845 85.835 ;
        RECT 129.325 83.500 129.605 89.860 ;
        RECT 130.175 83.500 130.475 90.320 ;
        RECT 131.315 82.755 131.615 89.910 ;
        RECT 133.600 88.615 133.975 96.900 ;
        RECT 135.345 87.895 135.645 98.890 ;
        RECT 136.490 86.780 136.870 97.035 ;
        RECT 137.360 84.625 137.795 98.200 ;
        RECT 193.065 97.400 193.580 107.450 ;
        RECT 194.750 96.045 195.335 106.825 ;
        RECT 196.590 104.390 196.945 118.180 ;
        RECT 259.935 117.550 260.385 128.050 ;
        RECT 198.215 105.245 198.575 116.580 ;
        RECT 261.100 116.010 261.585 125.250 ;
        RECT 267.515 115.765 267.920 127.295 ;
        RECT 269.590 117.665 269.980 128.765 ;
        RECT 272.995 121.255 273.350 132.340 ;
        RECT 276.740 130.980 277.030 133.040 ;
        RECT 279.510 131.580 280.010 134.630 ;
        RECT 284.480 131.490 284.890 134.585 ;
        RECT 283.520 129.830 283.830 129.860 ;
        RECT 274.320 126.110 274.790 129.100 ;
        RECT 276.670 123.125 276.985 125.495 ;
        RECT 278.290 125.170 278.710 129.135 ;
        RECT 274.955 120.415 275.335 121.790 ;
        RECT 277.395 119.385 277.740 121.845 ;
        RECT 279.030 121.065 279.355 123.830 ;
        RECT 280.015 123.100 280.420 126.430 ;
        RECT 283.520 123.730 283.835 129.830 ;
        RECT 284.665 120.125 285.035 129.225 ;
        RECT 285.610 121.190 285.900 133.025 ;
        RECT 289.060 131.465 289.470 134.560 ;
        RECT 293.515 130.920 293.825 133.435 ;
        RECT 297.765 132.620 298.145 133.000 ;
        RECT 299.895 132.620 300.275 133.000 ;
        RECT 286.505 123.685 286.835 129.880 ;
        RECT 289.410 123.155 289.865 126.430 ;
        RECT 291.770 125.170 292.315 129.110 ;
        RECT 295.825 126.110 296.260 129.120 ;
        RECT 290.965 121.065 291.290 123.830 ;
        RECT 293.480 123.160 293.895 125.550 ;
        RECT 297.020 121.735 297.350 132.430 ;
        RECT 298.455 126.070 298.840 131.855 ;
        RECT 295.210 120.330 295.545 121.680 ;
        RECT 298.815 121.315 299.240 125.590 ;
        RECT 300.515 123.080 300.815 130.120 ;
        RECT 301.635 122.475 301.935 129.405 ;
        RECT 302.945 123.075 303.245 129.425 ;
        RECT 297.475 120.405 297.855 120.785 ;
        RECT 299.670 120.390 300.050 120.770 ;
        RECT 303.540 120.330 303.830 130.110 ;
        RECT 304.260 123.105 304.555 129.930 ;
        RECT 305.390 122.565 305.690 129.375 ;
        RECT 306.180 123.160 306.490 133.200 ;
        RECT 315.370 131.445 315.750 131.825 ;
        RECT 306.975 123.090 307.275 129.920 ;
        RECT 308.100 122.475 308.400 129.415 ;
        RECT 309.550 122.350 309.830 125.385 ;
        RECT 310.310 123.050 310.590 129.410 ;
        RECT 311.160 123.050 311.460 129.870 ;
        RECT 312.300 122.305 312.600 129.460 ;
        RECT 312.945 126.495 313.325 126.875 ;
        RECT 312.945 124.440 313.325 124.820 ;
        RECT 314.795 124.320 315.110 128.645 ;
        RECT 315.405 126.395 315.685 127.925 ;
        RECT 315.975 123.080 316.275 130.120 ;
        RECT 317.095 122.475 317.395 129.405 ;
        RECT 317.750 123.835 318.050 127.895 ;
        RECT 318.405 123.075 318.705 129.425 ;
        RECT 315.270 121.270 315.650 121.650 ;
        RECT 319.000 120.865 319.290 130.110 ;
        RECT 319.720 123.105 320.015 129.930 ;
        RECT 320.850 122.565 321.150 129.375 ;
        RECT 321.640 123.160 321.950 131.895 ;
        RECT 322.435 123.090 322.735 129.920 ;
        RECT 323.560 122.475 323.860 129.415 ;
        RECT 324.240 123.820 324.520 127.910 ;
        RECT 325.010 122.350 325.290 125.385 ;
        RECT 325.770 123.050 326.050 129.410 ;
        RECT 326.620 123.050 326.920 129.870 ;
        RECT 327.760 122.305 328.060 129.460 ;
        RECT 329.945 128.095 330.320 136.295 ;
        RECT 331.690 127.290 331.990 138.285 ;
        RECT 332.880 126.290 333.260 136.545 ;
        RECT 333.750 124.135 334.185 137.710 ;
        RECT 389.455 136.910 389.970 146.960 ;
        RECT 391.140 135.555 391.725 146.335 ;
        RECT 392.780 143.880 393.135 157.670 ;
        RECT 456.125 157.040 456.575 167.305 ;
        RECT 394.405 144.735 394.765 156.070 ;
        RECT 457.290 155.500 457.775 164.385 ;
        RECT 463.595 155.125 464.000 166.655 ;
        RECT 465.670 157.025 466.060 168.125 ;
        RECT 469.440 160.575 469.795 171.660 ;
        RECT 473.185 170.300 473.475 172.360 ;
        RECT 475.955 170.900 476.455 173.950 ;
        RECT 480.925 170.810 481.335 173.905 ;
        RECT 479.965 169.150 480.275 169.180 ;
        RECT 470.765 165.430 471.235 168.420 ;
        RECT 473.115 162.445 473.430 164.815 ;
        RECT 474.735 164.490 475.155 168.455 ;
        RECT 471.400 159.735 471.780 161.110 ;
        RECT 473.840 158.705 474.185 161.165 ;
        RECT 475.475 160.385 475.800 163.150 ;
        RECT 476.460 162.420 476.865 165.750 ;
        RECT 479.965 163.050 480.280 169.150 ;
        RECT 481.110 159.445 481.480 168.545 ;
        RECT 482.055 160.510 482.345 172.345 ;
        RECT 485.505 170.785 485.915 173.880 ;
        RECT 489.960 170.240 490.270 172.755 ;
        RECT 494.210 171.940 494.590 172.320 ;
        RECT 496.340 171.940 496.720 172.320 ;
        RECT 482.950 163.005 483.280 169.200 ;
        RECT 485.855 162.475 486.310 165.750 ;
        RECT 488.215 164.490 488.760 168.430 ;
        RECT 492.270 165.430 492.705 168.440 ;
        RECT 487.410 160.385 487.735 163.150 ;
        RECT 489.925 162.480 490.340 164.870 ;
        RECT 493.465 161.055 493.795 171.750 ;
        RECT 494.900 165.390 495.285 171.175 ;
        RECT 491.655 159.650 491.990 161.000 ;
        RECT 495.260 160.635 495.685 164.910 ;
        RECT 496.960 162.400 497.260 169.440 ;
        RECT 498.080 161.795 498.380 168.725 ;
        RECT 499.390 162.395 499.690 168.745 ;
        RECT 493.920 159.725 494.300 160.105 ;
        RECT 496.115 159.710 496.495 160.090 ;
        RECT 499.985 159.650 500.275 169.430 ;
        RECT 500.705 162.425 501.000 169.250 ;
        RECT 501.835 161.885 502.135 168.695 ;
        RECT 502.625 162.480 502.935 172.520 ;
        RECT 511.815 170.765 512.195 171.145 ;
        RECT 503.420 162.410 503.720 169.240 ;
        RECT 504.545 161.795 504.845 168.735 ;
        RECT 505.995 161.670 506.275 164.705 ;
        RECT 506.755 162.370 507.035 168.730 ;
        RECT 507.605 162.370 507.905 169.190 ;
        RECT 508.745 161.625 509.045 168.780 ;
        RECT 509.390 165.815 509.770 166.195 ;
        RECT 509.390 163.760 509.770 164.140 ;
        RECT 511.240 163.640 511.555 167.965 ;
        RECT 511.850 165.715 512.130 167.245 ;
        RECT 512.420 162.400 512.720 169.440 ;
        RECT 514.195 163.155 514.495 167.215 ;
        RECT 511.715 160.590 512.095 160.970 ;
        RECT 515.445 160.185 515.735 169.430 ;
        RECT 517.295 161.885 517.595 168.695 ;
        RECT 518.085 162.480 518.395 171.215 ;
        RECT 518.880 162.410 519.180 169.240 ;
        RECT 520.685 163.140 520.965 167.230 ;
        RECT 521.455 161.670 521.735 164.705 ;
        RECT 524.205 161.625 524.505 168.780 ;
        RECT 561.045 160.700 561.360 171.750 ;
        RECT 564.880 171.045 565.280 174.095 ;
        RECT 569.800 170.955 570.210 174.050 ;
        RECT 574.380 170.930 574.790 174.025 ;
        RECT 562.715 158.850 563.060 161.310 ;
        RECT 579.830 161.185 580.145 171.870 ;
        RECT 585.015 163.975 585.465 168.135 ;
        RECT 594.475 167.670 594.855 168.050 ;
        RECT 586.715 166.955 587.240 167.395 ;
        RECT 594.465 166.920 594.845 167.300 ;
        RECT 398.055 147.945 398.435 148.325 ;
        RECT 398.045 147.195 398.425 147.575 ;
        RECT 398.090 146.510 398.470 146.890 ;
        RECT 398.055 145.840 398.435 146.220 ;
        RECT 398.770 142.765 399.070 149.805 ;
        RECT 399.890 142.160 400.190 149.090 ;
        RECT 400.545 143.520 400.845 147.580 ;
        RECT 401.200 142.760 401.500 149.110 ;
        RECT 401.795 144.635 402.115 149.795 ;
        RECT 402.515 142.790 402.810 149.615 ;
        RECT 403.645 142.250 403.945 149.060 ;
        RECT 404.435 142.845 404.745 149.035 ;
        RECT 405.230 142.775 405.530 149.605 ;
        RECT 406.355 142.160 406.655 149.100 ;
        RECT 407.035 143.505 407.315 147.595 ;
        RECT 407.805 142.035 408.085 145.070 ;
        RECT 408.565 142.735 408.870 149.095 ;
        RECT 409.415 142.735 409.715 149.555 ;
        RECT 410.555 141.990 410.855 149.145 ;
        RECT 411.220 147.945 411.600 148.325 ;
        RECT 413.490 147.945 413.870 148.350 ;
        RECT 411.225 147.195 411.605 147.575 ;
        RECT 413.495 147.195 413.875 147.600 ;
        RECT 411.225 146.180 411.605 146.560 ;
        RECT 413.010 144.760 413.330 146.890 ;
        RECT 411.440 141.470 411.820 144.490 ;
        RECT 413.620 143.920 413.900 146.325 ;
        RECT 414.230 142.765 414.530 149.805 ;
        RECT 415.350 142.160 415.650 149.090 ;
        RECT 416.005 143.520 416.305 147.580 ;
        RECT 416.660 142.760 416.960 149.110 ;
        RECT 417.255 144.635 417.580 149.795 ;
        RECT 417.975 142.790 418.270 149.615 ;
        RECT 419.105 142.250 419.405 149.060 ;
        RECT 419.895 142.845 420.205 149.035 ;
        RECT 420.690 142.775 420.990 149.605 ;
        RECT 421.815 142.160 422.115 149.100 ;
        RECT 422.495 143.505 422.775 147.595 ;
        RECT 423.265 142.035 423.545 145.070 ;
        RECT 424.025 142.735 424.345 149.095 ;
        RECT 424.875 142.735 425.175 149.555 ;
        RECT 426.015 141.990 426.315 149.145 ;
        RECT 426.955 147.945 427.315 149.775 ;
        RECT 426.650 144.135 427.030 144.515 ;
        RECT 427.355 140.020 427.715 146.580 ;
        RECT 428.495 144.770 428.820 146.635 ;
        RECT 429.135 146.425 429.550 149.775 ;
        RECT 429.160 141.425 429.620 146.110 ;
        RECT 429.945 143.970 430.395 152.790 ;
        RECT 430.805 141.595 431.160 151.900 ;
        RECT 431.470 147.200 431.815 148.255 ;
        RECT 432.130 145.795 432.560 148.785 ;
        RECT 429.875 140.080 430.255 140.460 ;
        RECT 432.765 140.100 433.145 141.475 ;
        RECT 433.535 140.920 433.850 151.970 ;
        RECT 434.550 150.665 434.840 152.725 ;
        RECT 437.335 151.265 437.810 154.315 ;
        RECT 442.290 151.175 442.700 154.270 ;
        RECT 441.330 149.515 441.640 149.545 ;
        RECT 434.470 142.810 434.795 145.180 ;
        RECT 436.120 144.855 436.520 148.820 ;
        RECT 435.205 139.070 435.550 141.530 ;
        RECT 436.840 140.750 437.165 143.515 ;
        RECT 437.825 142.785 438.230 146.115 ;
        RECT 441.330 143.415 441.645 149.515 ;
        RECT 442.475 139.810 442.845 148.910 ;
        RECT 443.420 140.875 443.710 152.710 ;
        RECT 446.870 151.150 447.280 154.245 ;
        RECT 451.325 150.605 451.635 153.120 ;
        RECT 444.315 143.370 444.645 149.565 ;
        RECT 447.235 142.840 447.675 146.115 ;
        RECT 449.615 144.855 450.140 148.795 ;
        RECT 448.775 140.750 449.100 143.515 ;
        RECT 451.290 142.845 451.705 145.235 ;
        RECT 452.320 141.405 452.635 152.090 ;
        RECT 453.650 145.795 454.135 148.805 ;
        RECT 454.830 141.420 455.160 152.115 ;
        RECT 453.020 140.015 453.355 141.365 ;
        RECT 364.700 121.135 365.015 132.185 ;
        RECT 368.535 131.480 368.935 134.530 ;
        RECT 373.455 131.390 373.865 134.485 ;
        RECT 378.035 131.365 378.445 134.460 ;
        RECT 366.370 119.285 366.715 121.745 ;
        RECT 383.485 121.620 383.800 132.305 ;
        RECT 388.670 124.410 389.120 128.570 ;
        RECT 390.370 127.390 390.895 127.830 ;
        RECT 201.650 108.445 202.030 108.825 ;
        RECT 201.640 107.695 202.020 108.075 ;
        RECT 201.685 107.010 202.065 107.390 ;
        RECT 201.650 106.340 202.030 106.720 ;
        RECT 202.365 103.265 202.665 110.305 ;
        RECT 203.485 102.660 203.785 109.590 ;
        RECT 204.140 104.020 204.440 108.080 ;
        RECT 204.795 103.260 205.095 109.610 ;
        RECT 205.390 105.135 205.710 110.295 ;
        RECT 206.110 103.290 206.405 110.115 ;
        RECT 207.240 102.750 207.540 109.560 ;
        RECT 208.030 103.345 208.340 109.535 ;
        RECT 208.825 103.275 209.125 110.105 ;
        RECT 209.950 102.660 210.250 109.600 ;
        RECT 210.630 104.005 210.910 108.095 ;
        RECT 211.400 102.535 211.680 105.570 ;
        RECT 212.160 103.235 212.465 109.595 ;
        RECT 213.010 103.235 213.310 110.055 ;
        RECT 214.150 102.490 214.450 109.645 ;
        RECT 214.815 108.445 215.195 108.825 ;
        RECT 217.085 108.445 217.465 108.850 ;
        RECT 214.820 107.695 215.200 108.075 ;
        RECT 217.090 107.695 217.470 108.100 ;
        RECT 214.820 106.680 215.200 107.060 ;
        RECT 216.605 105.260 216.925 107.390 ;
        RECT 215.035 101.970 215.415 104.990 ;
        RECT 217.215 104.420 217.495 106.825 ;
        RECT 217.825 103.265 218.125 110.305 ;
        RECT 218.945 102.660 219.245 109.590 ;
        RECT 219.600 104.020 219.900 108.080 ;
        RECT 220.255 103.260 220.555 109.610 ;
        RECT 220.850 105.135 221.175 110.295 ;
        RECT 221.570 103.290 221.865 110.115 ;
        RECT 222.700 102.750 223.000 109.560 ;
        RECT 223.490 103.345 223.800 109.535 ;
        RECT 224.285 103.275 224.585 110.105 ;
        RECT 225.410 102.660 225.710 109.600 ;
        RECT 226.090 104.005 226.370 108.095 ;
        RECT 226.860 102.535 227.140 105.570 ;
        RECT 227.620 103.235 227.940 109.595 ;
        RECT 228.470 103.235 228.770 110.055 ;
        RECT 229.610 102.490 229.910 109.645 ;
        RECT 230.550 108.445 230.910 110.275 ;
        RECT 230.245 104.635 230.625 105.015 ;
        RECT 230.950 100.520 231.310 107.080 ;
        RECT 232.090 105.270 232.415 107.135 ;
        RECT 232.730 106.925 233.145 110.275 ;
        RECT 232.755 101.925 233.215 106.610 ;
        RECT 233.540 104.470 233.990 113.290 ;
        RECT 234.400 102.095 234.755 112.400 ;
        RECT 235.065 107.700 235.410 108.755 ;
        RECT 235.725 106.295 236.155 109.285 ;
        RECT 233.470 100.580 233.850 100.960 ;
        RECT 236.360 100.600 236.740 101.975 ;
        RECT 237.130 101.420 237.445 112.470 ;
        RECT 238.145 111.165 238.435 113.225 ;
        RECT 240.930 111.765 241.405 114.815 ;
        RECT 245.885 111.675 246.295 114.770 ;
        RECT 244.925 110.015 245.235 110.045 ;
        RECT 238.065 103.310 238.390 105.680 ;
        RECT 239.715 105.355 240.115 109.320 ;
        RECT 238.800 99.570 239.145 102.030 ;
        RECT 240.435 101.250 240.760 104.015 ;
        RECT 241.420 103.285 241.825 106.615 ;
        RECT 244.925 103.915 245.240 110.015 ;
        RECT 246.070 100.310 246.440 109.410 ;
        RECT 247.015 101.375 247.305 113.210 ;
        RECT 250.465 111.650 250.875 114.745 ;
        RECT 254.920 111.105 255.230 113.620 ;
        RECT 247.910 103.870 248.240 110.065 ;
        RECT 250.830 103.340 251.270 106.615 ;
        RECT 253.210 105.355 253.735 109.295 ;
        RECT 252.370 101.250 252.695 104.015 ;
        RECT 254.885 103.345 255.300 105.735 ;
        RECT 255.915 101.905 256.230 112.590 ;
        RECT 257.245 106.295 257.730 109.305 ;
        RECT 258.425 101.920 258.755 112.615 ;
        RECT 256.615 100.515 256.950 101.865 ;
        RECT 168.270 81.680 168.585 92.730 ;
        RECT 172.105 92.025 172.505 95.075 ;
        RECT 177.025 91.935 177.435 95.030 ;
        RECT 181.605 91.910 182.015 95.005 ;
        RECT 169.940 79.830 170.285 82.290 ;
        RECT 187.055 82.165 187.370 92.850 ;
        RECT 192.240 84.955 192.690 89.115 ;
        RECT 193.940 87.935 194.465 88.375 ;
        RECT 5.285 68.975 5.665 69.355 ;
        RECT 5.275 68.225 5.655 68.605 ;
        RECT 5.320 67.540 5.700 67.920 ;
        RECT 5.285 66.870 5.665 67.250 ;
        RECT 6.000 63.795 6.300 70.835 ;
        RECT 7.120 63.190 7.420 70.120 ;
        RECT 7.775 64.550 8.075 68.610 ;
        RECT 8.430 63.790 8.730 70.140 ;
        RECT 9.025 65.665 9.345 70.825 ;
        RECT 9.745 63.820 10.040 70.645 ;
        RECT 10.875 63.280 11.175 70.090 ;
        RECT 11.665 63.875 11.975 70.065 ;
        RECT 12.460 63.805 12.760 70.635 ;
        RECT 13.585 63.190 13.885 70.130 ;
        RECT 14.265 64.535 14.545 68.625 ;
        RECT 15.035 63.065 15.315 66.100 ;
        RECT 15.795 63.765 16.100 70.125 ;
        RECT 16.645 63.765 16.945 70.585 ;
        RECT 17.785 63.020 18.085 70.175 ;
        RECT 18.450 68.975 18.830 69.355 ;
        RECT 20.720 68.975 21.100 69.380 ;
        RECT 18.455 68.225 18.835 68.605 ;
        RECT 20.725 68.225 21.105 68.630 ;
        RECT 18.455 67.210 18.835 67.590 ;
        RECT 20.240 65.790 20.560 67.920 ;
        RECT 18.670 62.500 19.050 65.520 ;
        RECT 20.850 64.950 21.130 67.355 ;
        RECT 21.460 63.795 21.760 70.835 ;
        RECT 22.580 63.190 22.880 70.120 ;
        RECT 23.235 64.550 23.535 68.610 ;
        RECT 23.890 63.790 24.190 70.140 ;
        RECT 24.485 65.665 24.810 70.825 ;
        RECT 25.205 63.820 25.500 70.645 ;
        RECT 26.335 63.280 26.635 70.090 ;
        RECT 27.125 63.875 27.435 70.065 ;
        RECT 27.920 63.805 28.220 70.635 ;
        RECT 29.045 63.190 29.345 70.130 ;
        RECT 29.725 64.535 30.005 68.625 ;
        RECT 30.495 63.065 30.775 66.100 ;
        RECT 31.255 63.765 31.575 70.125 ;
        RECT 32.105 63.765 32.405 70.585 ;
        RECT 33.245 63.020 33.545 70.175 ;
        RECT 34.185 68.975 34.545 70.805 ;
        RECT 33.880 65.165 34.260 65.545 ;
        RECT 34.585 61.050 34.945 67.610 ;
        RECT 35.725 65.800 36.050 67.665 ;
        RECT 36.365 67.455 36.780 70.805 ;
        RECT 36.390 62.455 36.850 67.140 ;
        RECT 37.175 65.000 37.625 73.820 ;
        RECT 38.035 62.625 38.390 72.930 ;
        RECT 38.700 68.230 39.045 69.285 ;
        RECT 39.360 66.825 39.790 69.815 ;
        RECT 37.105 61.110 37.485 61.490 ;
        RECT 39.995 61.130 40.375 62.505 ;
        RECT 40.765 61.950 41.080 73.000 ;
        RECT 41.780 71.695 42.070 73.755 ;
        RECT 44.565 72.295 45.040 75.345 ;
        RECT 49.520 72.205 49.930 75.300 ;
        RECT 48.560 70.545 48.870 70.575 ;
        RECT 41.700 63.840 42.025 66.210 ;
        RECT 43.350 65.885 43.750 69.850 ;
        RECT 42.435 60.100 42.780 62.560 ;
        RECT 44.070 61.780 44.395 64.545 ;
        RECT 45.055 63.815 45.460 67.145 ;
        RECT 48.560 64.445 48.875 70.545 ;
        RECT 49.705 60.840 50.075 69.940 ;
        RECT 50.650 61.905 50.940 73.740 ;
        RECT 54.100 72.180 54.510 75.275 ;
        RECT 58.555 71.635 58.865 74.150 ;
        RECT 51.545 64.400 51.875 70.595 ;
        RECT 54.465 63.870 54.905 67.145 ;
        RECT 56.845 65.885 57.370 69.825 ;
        RECT 56.005 61.780 56.330 64.545 ;
        RECT 58.520 63.875 58.935 66.265 ;
        RECT 59.550 62.435 59.865 73.120 ;
        RECT 60.880 66.825 61.365 69.835 ;
        RECT 62.060 62.450 62.390 73.145 ;
        RECT 60.250 61.045 60.585 62.395 ;
        RECT -78.225 42.040 -77.910 53.090 ;
        RECT -74.390 52.385 -73.990 55.435 ;
        RECT -69.470 52.295 -69.060 55.390 ;
        RECT -64.890 52.270 -64.480 55.365 ;
        RECT -76.555 40.190 -76.210 42.650 ;
        RECT -59.440 42.525 -59.125 53.210 ;
        RECT -55.750 45.320 -55.335 48.135 ;
        RECT -55.010 46.905 -54.625 48.800 ;
        RECT -27.900 42.120 -27.585 53.170 ;
        RECT -24.065 52.465 -23.665 55.515 ;
        RECT -19.145 52.375 -18.735 55.470 ;
        RECT -14.565 52.350 -14.155 55.445 ;
        RECT -26.230 40.270 -25.885 42.730 ;
        RECT -9.115 42.605 -8.800 53.290 ;
        RECT -3.930 45.395 -3.480 49.555 ;
        RECT -2.230 48.375 -1.705 48.815 ;
        RECT -0.030 45.075 0.325 58.985 ;
        RECT 63.315 58.355 63.765 68.620 ;
        RECT 1.595 45.995 1.955 57.385 ;
        RECT 64.480 56.815 64.965 65.700 ;
        RECT 71.310 56.170 71.715 68.050 ;
        RECT 73.385 58.070 73.775 69.650 ;
        RECT 76.655 61.990 77.010 73.075 ;
        RECT 80.400 71.715 80.690 73.775 ;
        RECT 83.170 72.315 83.670 75.365 ;
        RECT 88.140 72.225 88.550 75.320 ;
        RECT 87.180 70.565 87.490 70.595 ;
        RECT 77.980 66.845 78.450 69.835 ;
        RECT 80.330 63.860 80.645 66.230 ;
        RECT 81.950 65.905 82.370 69.870 ;
        RECT 78.615 61.150 78.995 62.525 ;
        RECT 81.055 60.120 81.400 62.580 ;
        RECT 82.690 61.800 83.015 64.565 ;
        RECT 83.675 63.835 84.080 67.165 ;
        RECT 87.180 64.465 87.495 70.565 ;
        RECT 88.325 60.860 88.695 69.960 ;
        RECT 89.270 61.925 89.560 73.760 ;
        RECT 92.720 72.200 93.130 75.295 ;
        RECT 97.175 71.655 97.485 74.170 ;
        RECT 101.425 73.355 101.805 73.735 ;
        RECT 103.555 73.355 103.935 73.735 ;
        RECT 90.165 64.420 90.495 70.615 ;
        RECT 93.070 63.890 93.525 67.165 ;
        RECT 95.430 65.905 95.975 69.845 ;
        RECT 99.485 66.845 99.920 69.855 ;
        RECT 94.625 61.800 94.950 64.565 ;
        RECT 97.140 63.895 97.555 66.285 ;
        RECT 100.680 62.470 101.010 73.165 ;
        RECT 102.115 66.805 102.500 72.590 ;
        RECT 98.870 61.065 99.205 62.415 ;
        RECT 102.475 62.050 102.900 66.325 ;
        RECT 104.175 63.815 104.475 70.855 ;
        RECT 105.295 63.210 105.595 70.140 ;
        RECT 106.605 63.810 106.905 70.160 ;
        RECT 101.135 61.140 101.515 61.520 ;
        RECT 103.330 61.125 103.710 61.505 ;
        RECT 107.200 61.065 107.490 70.845 ;
        RECT 107.920 63.840 108.215 70.665 ;
        RECT 109.050 63.300 109.350 70.110 ;
        RECT 109.840 63.895 110.150 73.935 ;
        RECT 119.030 72.180 119.410 72.560 ;
        RECT 110.635 63.825 110.935 70.655 ;
        RECT 111.760 63.210 112.060 70.150 ;
        RECT 113.210 63.085 113.490 66.120 ;
        RECT 113.970 63.785 114.250 70.145 ;
        RECT 114.820 63.785 115.120 70.605 ;
        RECT 115.960 63.040 116.260 70.195 ;
        RECT 116.605 67.230 116.985 67.610 ;
        RECT 116.605 65.175 116.985 65.555 ;
        RECT 118.455 65.055 118.770 69.380 ;
        RECT 119.065 67.130 119.345 68.660 ;
        RECT 119.635 63.815 119.935 70.855 ;
        RECT 120.755 63.210 121.055 70.140 ;
        RECT 121.410 64.570 121.710 68.630 ;
        RECT 122.065 63.810 122.365 70.160 ;
        RECT 118.930 62.005 119.310 62.385 ;
        RECT 122.660 61.600 122.950 70.845 ;
        RECT 123.380 63.840 123.675 70.665 ;
        RECT 124.510 63.300 124.810 70.110 ;
        RECT 125.300 63.895 125.610 72.630 ;
        RECT 126.095 63.825 126.395 70.655 ;
        RECT 127.220 63.210 127.520 70.150 ;
        RECT 127.900 64.555 128.180 68.645 ;
        RECT 128.670 63.085 128.950 66.120 ;
        RECT 129.430 63.785 129.710 70.145 ;
        RECT 130.280 63.785 130.580 70.605 ;
        RECT 131.420 63.040 131.720 70.195 ;
        RECT 133.500 68.915 133.875 77.195 ;
        RECT 135.245 68.075 135.545 79.185 ;
        RECT 136.490 67.070 136.870 77.325 ;
        RECT 137.360 64.915 137.795 78.490 ;
        RECT 193.070 77.690 193.585 87.740 ;
        RECT 194.755 76.335 195.340 87.115 ;
        RECT 196.545 84.600 196.900 98.390 ;
        RECT 259.890 97.760 260.340 108.250 ;
        RECT 198.170 85.505 198.530 96.790 ;
        RECT 261.055 96.220 261.540 105.380 ;
        RECT 267.515 96.030 267.920 107.560 ;
        RECT 269.590 97.930 269.980 109.030 ;
        RECT 272.995 101.460 273.350 112.545 ;
        RECT 276.740 111.185 277.030 113.245 ;
        RECT 279.510 111.785 280.010 114.835 ;
        RECT 284.480 111.695 284.890 114.790 ;
        RECT 283.520 110.035 283.830 110.065 ;
        RECT 274.320 106.315 274.790 109.305 ;
        RECT 276.670 103.330 276.985 105.700 ;
        RECT 278.290 105.375 278.710 109.340 ;
        RECT 274.955 100.620 275.335 101.995 ;
        RECT 277.395 99.590 277.740 102.050 ;
        RECT 279.030 101.270 279.355 104.035 ;
        RECT 280.015 103.305 280.420 106.635 ;
        RECT 283.520 103.935 283.835 110.035 ;
        RECT 284.665 100.330 285.035 109.430 ;
        RECT 285.610 101.395 285.900 113.230 ;
        RECT 289.060 111.670 289.470 114.765 ;
        RECT 293.515 111.125 293.825 113.640 ;
        RECT 297.765 112.825 298.145 113.205 ;
        RECT 299.895 112.825 300.275 113.205 ;
        RECT 286.505 103.890 286.835 110.085 ;
        RECT 289.410 103.360 289.865 106.635 ;
        RECT 291.770 105.375 292.315 109.315 ;
        RECT 295.825 106.315 296.260 109.325 ;
        RECT 290.965 101.270 291.290 104.035 ;
        RECT 293.480 103.365 293.895 105.755 ;
        RECT 297.020 101.940 297.350 112.635 ;
        RECT 298.455 106.275 298.840 112.060 ;
        RECT 295.210 100.535 295.545 101.885 ;
        RECT 298.815 101.520 299.240 105.795 ;
        RECT 300.515 103.285 300.815 110.325 ;
        RECT 301.635 102.680 301.935 109.610 ;
        RECT 302.945 103.280 303.245 109.630 ;
        RECT 297.475 100.610 297.855 100.990 ;
        RECT 299.670 100.595 300.050 100.975 ;
        RECT 303.540 100.535 303.830 110.315 ;
        RECT 304.260 103.310 304.555 110.135 ;
        RECT 305.390 102.770 305.690 109.580 ;
        RECT 306.180 103.365 306.490 113.405 ;
        RECT 315.370 111.650 315.750 112.030 ;
        RECT 306.975 103.295 307.275 110.125 ;
        RECT 308.100 102.680 308.400 109.620 ;
        RECT 309.550 102.555 309.830 105.590 ;
        RECT 310.310 103.255 310.590 109.615 ;
        RECT 311.160 103.255 311.460 110.075 ;
        RECT 312.300 102.510 312.600 109.665 ;
        RECT 312.945 106.700 313.325 107.080 ;
        RECT 312.945 104.645 313.325 105.025 ;
        RECT 314.795 104.525 315.110 108.850 ;
        RECT 315.405 106.600 315.685 108.130 ;
        RECT 315.975 103.285 316.275 110.325 ;
        RECT 317.095 102.680 317.395 109.610 ;
        RECT 317.750 104.040 318.050 108.100 ;
        RECT 318.405 103.280 318.705 109.630 ;
        RECT 315.270 101.475 315.650 101.855 ;
        RECT 319.000 101.070 319.290 110.315 ;
        RECT 319.720 103.310 320.015 110.135 ;
        RECT 320.850 102.770 321.150 109.580 ;
        RECT 321.640 103.365 321.950 112.100 ;
        RECT 322.435 103.295 322.735 110.125 ;
        RECT 323.560 102.680 323.860 109.620 ;
        RECT 324.240 104.025 324.520 108.115 ;
        RECT 325.010 102.555 325.290 105.590 ;
        RECT 325.770 103.255 326.050 109.615 ;
        RECT 326.620 103.255 326.920 110.075 ;
        RECT 327.760 102.510 328.060 109.665 ;
        RECT 329.965 108.435 330.340 116.635 ;
        RECT 331.710 107.630 332.010 118.625 ;
        RECT 332.880 106.495 333.260 116.750 ;
        RECT 333.750 104.340 334.185 117.915 ;
        RECT 389.605 117.195 390.120 127.245 ;
        RECT 391.290 115.840 391.875 126.620 ;
        RECT 392.780 124.115 393.135 138.170 ;
        RECT 456.125 137.540 456.575 147.655 ;
        RECT 394.405 124.920 394.765 136.570 ;
        RECT 457.290 136.000 457.775 144.755 ;
        RECT 463.895 135.375 464.300 146.905 ;
        RECT 465.970 137.275 466.360 148.375 ;
        RECT 469.240 140.850 469.595 151.935 ;
        RECT 472.985 150.575 473.275 152.635 ;
        RECT 475.755 151.175 476.255 154.225 ;
        RECT 480.725 151.085 481.135 154.180 ;
        RECT 479.765 149.425 480.075 149.455 ;
        RECT 470.565 145.705 471.035 148.695 ;
        RECT 472.915 142.720 473.230 145.090 ;
        RECT 474.535 144.765 474.955 148.730 ;
        RECT 471.200 140.010 471.580 141.385 ;
        RECT 473.640 138.980 473.985 141.440 ;
        RECT 475.275 140.660 475.600 143.425 ;
        RECT 476.260 142.695 476.665 146.025 ;
        RECT 479.765 143.325 480.080 149.425 ;
        RECT 480.910 139.720 481.280 148.820 ;
        RECT 481.855 140.785 482.145 152.620 ;
        RECT 485.305 151.060 485.715 154.155 ;
        RECT 489.760 150.515 490.070 153.030 ;
        RECT 494.010 152.215 494.390 152.595 ;
        RECT 496.140 152.215 496.520 152.595 ;
        RECT 482.750 143.280 483.080 149.475 ;
        RECT 485.655 142.750 486.110 146.025 ;
        RECT 488.015 144.765 488.560 148.705 ;
        RECT 492.070 145.705 492.505 148.715 ;
        RECT 487.210 140.660 487.535 143.425 ;
        RECT 489.725 142.755 490.140 145.145 ;
        RECT 493.265 141.330 493.595 152.025 ;
        RECT 494.700 145.665 495.085 151.450 ;
        RECT 491.455 139.925 491.790 141.275 ;
        RECT 495.060 140.910 495.485 145.185 ;
        RECT 496.760 142.675 497.060 149.715 ;
        RECT 497.880 142.070 498.180 149.000 ;
        RECT 499.190 142.670 499.490 149.020 ;
        RECT 493.720 140.000 494.100 140.380 ;
        RECT 495.915 139.985 496.295 140.365 ;
        RECT 499.785 139.925 500.075 149.705 ;
        RECT 500.505 142.700 500.800 149.525 ;
        RECT 501.635 142.160 501.935 148.970 ;
        RECT 502.425 142.755 502.735 152.795 ;
        RECT 511.615 151.040 511.995 151.420 ;
        RECT 503.220 142.685 503.520 149.515 ;
        RECT 504.345 142.070 504.645 149.010 ;
        RECT 505.795 141.945 506.075 144.980 ;
        RECT 506.555 142.645 506.835 149.005 ;
        RECT 507.405 142.645 507.705 149.465 ;
        RECT 508.545 141.900 508.845 149.055 ;
        RECT 509.190 146.090 509.570 146.470 ;
        RECT 509.190 144.035 509.570 144.415 ;
        RECT 511.040 143.915 511.355 148.240 ;
        RECT 511.650 145.990 511.930 147.520 ;
        RECT 512.220 142.675 512.520 149.715 ;
        RECT 513.340 142.070 513.640 149.000 ;
        RECT 513.995 143.430 514.295 147.490 ;
        RECT 514.650 142.670 514.950 149.020 ;
        RECT 511.515 140.865 511.895 141.245 ;
        RECT 515.245 140.460 515.535 149.705 ;
        RECT 515.965 142.700 516.260 149.525 ;
        RECT 517.095 142.160 517.395 148.970 ;
        RECT 517.885 142.755 518.195 151.490 ;
        RECT 518.680 142.685 518.980 149.515 ;
        RECT 519.805 142.070 520.105 149.010 ;
        RECT 520.485 143.415 520.765 147.505 ;
        RECT 521.255 141.945 521.535 144.980 ;
        RECT 522.015 142.645 522.295 149.005 ;
        RECT 522.865 142.645 523.165 149.465 ;
        RECT 524.005 141.900 524.305 149.055 ;
        RECT 526.045 147.795 526.420 155.995 ;
        RECT 527.790 146.990 528.090 157.985 ;
        RECT 529.200 145.980 529.580 156.235 ;
        RECT 530.070 143.825 530.505 157.400 ;
        RECT 585.775 156.645 586.290 166.695 ;
        RECT 594.510 166.235 594.890 166.615 ;
        RECT 587.460 155.290 588.045 166.070 ;
        RECT 594.475 165.565 594.855 165.945 ;
        RECT 595.190 162.490 595.490 169.530 ;
        RECT 596.310 161.885 596.610 168.815 ;
        RECT 596.965 163.245 597.265 167.305 ;
        RECT 597.620 162.485 597.920 168.835 ;
        RECT 598.215 164.360 598.535 169.520 ;
        RECT 598.935 162.515 599.230 169.340 ;
        RECT 600.065 161.975 600.365 168.785 ;
        RECT 600.855 162.570 601.165 168.760 ;
        RECT 601.650 162.500 601.950 169.330 ;
        RECT 602.775 161.885 603.075 168.825 ;
        RECT 603.455 163.230 603.735 167.320 ;
        RECT 604.225 161.760 604.505 164.795 ;
        RECT 604.985 162.460 605.290 168.820 ;
        RECT 605.835 162.460 606.135 169.280 ;
        RECT 606.975 161.715 607.275 168.870 ;
        RECT 607.640 167.670 608.020 168.050 ;
        RECT 609.910 167.670 610.290 168.075 ;
        RECT 607.645 166.920 608.025 167.300 ;
        RECT 609.915 166.920 610.295 167.325 ;
        RECT 607.645 165.905 608.025 166.285 ;
        RECT 609.430 164.485 609.750 166.615 ;
        RECT 607.860 161.195 608.240 164.215 ;
        RECT 610.040 163.645 610.320 166.050 ;
        RECT 610.650 162.490 610.950 169.530 ;
        RECT 611.770 161.885 612.070 168.815 ;
        RECT 612.425 163.245 612.725 167.305 ;
        RECT 613.080 162.485 613.380 168.835 ;
        RECT 613.675 164.360 614.000 169.520 ;
        RECT 614.395 162.515 614.690 169.340 ;
        RECT 615.525 161.975 615.825 168.785 ;
        RECT 616.315 162.570 616.625 168.760 ;
        RECT 617.110 162.500 617.410 169.330 ;
        RECT 618.235 161.885 618.535 168.825 ;
        RECT 618.915 163.230 619.195 167.320 ;
        RECT 619.685 161.760 619.965 164.795 ;
        RECT 620.445 162.460 620.765 168.820 ;
        RECT 621.295 162.460 621.595 169.280 ;
        RECT 622.435 161.715 622.735 168.870 ;
        RECT 623.375 167.670 623.735 169.500 ;
        RECT 623.070 163.860 623.450 164.240 ;
        RECT 623.775 159.745 624.135 166.305 ;
        RECT 624.915 164.495 625.240 166.360 ;
        RECT 625.555 166.150 625.970 169.500 ;
        RECT 625.580 161.150 626.040 165.835 ;
        RECT 626.365 163.695 626.815 172.515 ;
        RECT 627.225 161.320 627.580 171.625 ;
        RECT 627.890 166.925 628.235 167.980 ;
        RECT 628.550 165.520 628.980 168.510 ;
        RECT 626.295 159.805 626.675 160.185 ;
        RECT 629.185 159.825 629.565 161.200 ;
        RECT 629.955 160.645 630.270 171.695 ;
        RECT 630.970 170.390 631.260 172.450 ;
        RECT 633.755 170.990 634.230 174.040 ;
        RECT 638.710 170.900 639.120 173.995 ;
        RECT 637.750 169.240 638.060 169.270 ;
        RECT 630.890 162.535 631.215 164.905 ;
        RECT 632.540 164.580 632.940 168.545 ;
        RECT 631.625 158.795 631.970 161.255 ;
        RECT 633.260 160.475 633.585 163.240 ;
        RECT 634.245 162.510 634.650 165.840 ;
        RECT 637.750 163.140 638.065 169.240 ;
        RECT 638.895 159.535 639.265 168.635 ;
        RECT 639.840 160.600 640.130 172.435 ;
        RECT 643.290 170.875 643.700 173.970 ;
        RECT 647.745 170.330 648.055 172.845 ;
        RECT 640.735 163.095 641.065 169.290 ;
        RECT 643.655 162.565 644.095 165.840 ;
        RECT 646.035 164.580 646.560 168.520 ;
        RECT 645.195 160.475 645.520 163.240 ;
        RECT 647.710 162.570 648.125 164.960 ;
        RECT 648.740 161.130 649.055 171.815 ;
        RECT 650.070 165.520 650.555 168.530 ;
        RECT 651.250 161.145 651.580 171.840 ;
        RECT 649.440 159.740 649.775 161.090 ;
        RECT 560.960 140.985 561.275 152.035 ;
        RECT 564.795 151.330 565.195 154.380 ;
        RECT 569.715 151.240 570.125 154.335 ;
        RECT 574.295 151.215 574.705 154.310 ;
        RECT 562.630 139.135 562.975 141.595 ;
        RECT 579.745 141.470 580.060 152.155 ;
        RECT 584.930 144.260 585.380 148.420 ;
        RECT 586.630 147.240 587.155 147.680 ;
        RECT 398.245 128.235 398.625 128.615 ;
        RECT 398.235 127.485 398.615 127.865 ;
        RECT 398.280 126.800 398.660 127.180 ;
        RECT 398.245 126.130 398.625 126.510 ;
        RECT 398.960 123.055 399.260 130.095 ;
        RECT 400.080 122.450 400.380 129.380 ;
        RECT 400.735 123.810 401.035 127.870 ;
        RECT 401.390 123.050 401.690 129.400 ;
        RECT 401.985 124.925 402.305 130.085 ;
        RECT 402.705 123.080 403.000 129.905 ;
        RECT 403.835 122.540 404.135 129.350 ;
        RECT 404.625 123.135 404.935 129.325 ;
        RECT 405.420 123.065 405.720 129.895 ;
        RECT 406.545 122.450 406.845 129.390 ;
        RECT 407.225 123.795 407.505 127.885 ;
        RECT 407.995 122.325 408.275 125.360 ;
        RECT 408.755 123.025 409.060 129.385 ;
        RECT 409.605 123.025 409.905 129.845 ;
        RECT 410.745 122.280 411.045 129.435 ;
        RECT 411.410 128.235 411.790 128.615 ;
        RECT 413.680 128.235 414.060 128.640 ;
        RECT 411.415 127.485 411.795 127.865 ;
        RECT 413.685 127.485 414.065 127.890 ;
        RECT 411.415 126.470 411.795 126.850 ;
        RECT 413.200 125.050 413.520 127.180 ;
        RECT 411.630 121.760 412.010 124.780 ;
        RECT 413.810 124.210 414.090 126.615 ;
        RECT 414.420 123.055 414.720 130.095 ;
        RECT 415.540 122.450 415.840 129.380 ;
        RECT 416.195 123.810 416.495 127.870 ;
        RECT 416.850 123.050 417.150 129.400 ;
        RECT 417.445 124.925 417.770 130.085 ;
        RECT 418.165 123.080 418.460 129.905 ;
        RECT 419.295 122.540 419.595 129.350 ;
        RECT 420.085 123.135 420.395 129.325 ;
        RECT 420.880 123.065 421.180 129.895 ;
        RECT 422.005 122.450 422.305 129.390 ;
        RECT 422.685 123.795 422.965 127.885 ;
        RECT 423.455 122.325 423.735 125.360 ;
        RECT 424.215 123.025 424.535 129.385 ;
        RECT 425.065 123.025 425.365 129.845 ;
        RECT 426.205 122.280 426.505 129.435 ;
        RECT 427.145 128.235 427.505 130.065 ;
        RECT 426.840 124.425 427.220 124.805 ;
        RECT 427.545 120.310 427.905 126.870 ;
        RECT 428.685 125.060 429.010 126.925 ;
        RECT 429.325 126.715 429.740 130.065 ;
        RECT 429.350 121.715 429.810 126.400 ;
        RECT 430.135 124.260 430.585 133.080 ;
        RECT 430.995 121.885 431.350 132.190 ;
        RECT 431.660 127.490 432.005 128.545 ;
        RECT 432.320 126.085 432.750 129.075 ;
        RECT 430.065 120.370 430.445 120.750 ;
        RECT 432.955 120.390 433.335 121.765 ;
        RECT 433.725 121.210 434.040 132.260 ;
        RECT 434.740 130.955 435.030 133.015 ;
        RECT 437.525 131.555 438.000 134.605 ;
        RECT 442.480 131.465 442.890 134.560 ;
        RECT 441.520 129.805 441.830 129.835 ;
        RECT 434.660 123.100 434.985 125.470 ;
        RECT 436.310 125.145 436.710 129.110 ;
        RECT 435.395 119.360 435.740 121.820 ;
        RECT 437.030 121.040 437.355 123.805 ;
        RECT 438.015 123.075 438.420 126.405 ;
        RECT 441.520 123.705 441.835 129.805 ;
        RECT 442.665 120.100 443.035 129.200 ;
        RECT 443.610 121.165 443.900 133.000 ;
        RECT 447.060 131.440 447.470 134.535 ;
        RECT 451.515 130.895 451.825 133.410 ;
        RECT 444.505 123.660 444.835 129.855 ;
        RECT 447.425 123.130 447.865 126.405 ;
        RECT 449.805 125.145 450.330 129.085 ;
        RECT 448.965 121.040 449.290 123.805 ;
        RECT 451.480 123.135 451.895 125.525 ;
        RECT 452.510 121.695 452.825 132.380 ;
        RECT 453.840 126.085 454.325 129.095 ;
        RECT 455.020 121.710 455.350 132.405 ;
        RECT 453.210 120.305 453.545 121.655 ;
        RECT 364.630 101.365 364.945 112.415 ;
        RECT 368.465 111.710 368.865 114.760 ;
        RECT 373.385 111.620 373.795 114.715 ;
        RECT 377.965 111.595 378.375 114.690 ;
        RECT 366.300 99.515 366.645 101.975 ;
        RECT 383.415 101.850 383.730 112.535 ;
        RECT 388.600 104.640 389.050 108.800 ;
        RECT 390.300 107.620 390.825 108.060 ;
        RECT 201.520 88.735 201.900 89.115 ;
        RECT 201.510 87.985 201.890 88.365 ;
        RECT 201.555 87.300 201.935 87.680 ;
        RECT 201.520 86.630 201.900 87.010 ;
        RECT 202.235 83.555 202.535 90.595 ;
        RECT 203.355 82.950 203.655 89.880 ;
        RECT 204.010 84.310 204.310 88.370 ;
        RECT 204.665 83.550 204.965 89.900 ;
        RECT 205.260 85.425 205.580 90.585 ;
        RECT 205.980 83.580 206.275 90.405 ;
        RECT 207.110 83.040 207.410 89.850 ;
        RECT 207.900 83.635 208.210 89.825 ;
        RECT 208.695 83.565 208.995 90.395 ;
        RECT 209.820 82.950 210.120 89.890 ;
        RECT 210.500 84.295 210.780 88.385 ;
        RECT 211.270 82.825 211.550 85.860 ;
        RECT 212.030 83.525 212.335 89.885 ;
        RECT 212.880 83.525 213.180 90.345 ;
        RECT 214.020 82.780 214.320 89.935 ;
        RECT 214.685 88.735 215.065 89.115 ;
        RECT 216.955 88.735 217.335 89.140 ;
        RECT 214.690 87.985 215.070 88.365 ;
        RECT 216.960 87.985 217.340 88.390 ;
        RECT 214.690 86.970 215.070 87.350 ;
        RECT 216.475 85.550 216.795 87.680 ;
        RECT 214.905 82.260 215.285 85.280 ;
        RECT 217.085 84.710 217.365 87.115 ;
        RECT 217.695 83.555 217.995 90.595 ;
        RECT 218.815 82.950 219.115 89.880 ;
        RECT 219.470 84.310 219.770 88.370 ;
        RECT 220.125 83.550 220.425 89.900 ;
        RECT 220.720 85.425 221.045 90.585 ;
        RECT 221.440 83.580 221.735 90.405 ;
        RECT 222.570 83.040 222.870 89.850 ;
        RECT 223.360 83.635 223.670 89.825 ;
        RECT 224.155 83.565 224.455 90.395 ;
        RECT 225.280 82.950 225.580 89.890 ;
        RECT 225.960 84.295 226.240 88.385 ;
        RECT 226.730 82.825 227.010 85.860 ;
        RECT 227.490 83.525 227.810 89.885 ;
        RECT 228.340 83.525 228.640 90.345 ;
        RECT 229.480 82.780 229.780 89.935 ;
        RECT 230.420 88.735 230.780 90.565 ;
        RECT 230.115 84.925 230.495 85.305 ;
        RECT 230.820 80.810 231.180 87.370 ;
        RECT 231.960 85.560 232.285 87.425 ;
        RECT 232.600 87.215 233.015 90.565 ;
        RECT 232.625 82.215 233.085 86.900 ;
        RECT 233.410 84.760 233.860 93.580 ;
        RECT 234.270 82.385 234.625 92.690 ;
        RECT 234.935 87.990 235.280 89.045 ;
        RECT 235.595 86.585 236.025 89.575 ;
        RECT 233.340 80.870 233.720 81.250 ;
        RECT 236.230 80.890 236.610 82.265 ;
        RECT 237.000 81.710 237.315 92.760 ;
        RECT 238.015 91.455 238.305 93.515 ;
        RECT 240.800 92.055 241.275 95.105 ;
        RECT 245.755 91.965 246.165 95.060 ;
        RECT 244.795 90.305 245.105 90.335 ;
        RECT 237.935 83.600 238.260 85.970 ;
        RECT 239.585 85.645 239.985 89.610 ;
        RECT 238.670 79.860 239.015 82.320 ;
        RECT 240.305 81.540 240.630 84.305 ;
        RECT 241.290 83.575 241.695 86.905 ;
        RECT 244.795 84.205 245.110 90.305 ;
        RECT 245.940 80.600 246.310 89.700 ;
        RECT 246.885 81.665 247.175 93.500 ;
        RECT 250.335 91.940 250.745 95.035 ;
        RECT 254.790 91.395 255.100 93.910 ;
        RECT 247.780 84.160 248.110 90.355 ;
        RECT 250.700 83.630 251.140 86.905 ;
        RECT 253.080 85.645 253.605 89.585 ;
        RECT 252.240 81.540 252.565 84.305 ;
        RECT 254.755 83.635 255.170 86.025 ;
        RECT 255.785 82.195 256.100 92.880 ;
        RECT 257.115 86.585 257.600 89.595 ;
        RECT 258.295 82.210 258.625 92.905 ;
        RECT 256.485 80.805 256.820 82.155 ;
        RECT 168.200 61.850 168.515 72.900 ;
        RECT 172.035 72.195 172.435 75.245 ;
        RECT 176.955 72.105 177.365 75.200 ;
        RECT 181.535 72.080 181.945 75.175 ;
        RECT 169.870 60.000 170.215 62.460 ;
        RECT 186.985 62.335 187.300 73.020 ;
        RECT 192.170 65.125 192.620 69.285 ;
        RECT 193.870 68.105 194.395 68.545 ;
        RECT 5.235 49.165 5.615 49.545 ;
        RECT 5.225 48.415 5.605 48.795 ;
        RECT 5.270 47.730 5.650 48.110 ;
        RECT 5.235 47.060 5.615 47.440 ;
        RECT 5.950 43.985 6.250 51.025 ;
        RECT 7.070 43.380 7.370 50.310 ;
        RECT 7.725 44.740 8.025 48.800 ;
        RECT 8.380 43.980 8.680 50.330 ;
        RECT 8.975 45.855 9.295 51.015 ;
        RECT 9.695 44.010 9.990 50.835 ;
        RECT 10.825 43.470 11.125 50.280 ;
        RECT 11.615 44.065 11.925 50.255 ;
        RECT 12.410 43.995 12.710 50.825 ;
        RECT 13.535 43.380 13.835 50.320 ;
        RECT 14.215 44.725 14.495 48.815 ;
        RECT 14.985 43.255 15.265 46.290 ;
        RECT 15.745 43.955 16.050 50.315 ;
        RECT 16.595 43.955 16.895 50.775 ;
        RECT 17.735 43.210 18.035 50.365 ;
        RECT 18.400 49.165 18.780 49.545 ;
        RECT 20.670 49.165 21.050 49.570 ;
        RECT 18.405 48.415 18.785 48.795 ;
        RECT 20.675 48.415 21.055 48.820 ;
        RECT 18.405 47.400 18.785 47.780 ;
        RECT 20.190 45.980 20.510 48.110 ;
        RECT 18.620 42.690 19.000 45.710 ;
        RECT 20.800 45.140 21.080 47.545 ;
        RECT 21.410 43.985 21.710 51.025 ;
        RECT 22.530 43.380 22.830 50.310 ;
        RECT 23.185 44.740 23.485 48.800 ;
        RECT 23.840 43.980 24.140 50.330 ;
        RECT 24.435 45.855 24.760 51.015 ;
        RECT 25.155 44.010 25.450 50.835 ;
        RECT 26.285 43.470 26.585 50.280 ;
        RECT 27.075 44.065 27.385 50.255 ;
        RECT 27.870 43.995 28.170 50.825 ;
        RECT 28.995 43.380 29.295 50.320 ;
        RECT 29.675 44.725 29.955 48.815 ;
        RECT 30.445 43.255 30.725 46.290 ;
        RECT 31.205 43.955 31.525 50.315 ;
        RECT 32.055 43.955 32.355 50.775 ;
        RECT 33.195 43.210 33.495 50.365 ;
        RECT 34.135 49.165 34.495 50.995 ;
        RECT 33.830 45.355 34.210 45.735 ;
        RECT 34.535 41.240 34.895 47.800 ;
        RECT 35.675 45.990 36.000 47.855 ;
        RECT 36.315 47.645 36.730 50.995 ;
        RECT 36.340 42.645 36.800 47.330 ;
        RECT 37.125 45.190 37.575 54.010 ;
        RECT 37.985 42.815 38.340 53.120 ;
        RECT 38.650 48.420 38.995 49.475 ;
        RECT 39.310 47.015 39.740 50.005 ;
        RECT 37.055 41.300 37.435 41.680 ;
        RECT 39.945 41.320 40.325 42.695 ;
        RECT 40.715 42.140 41.030 53.190 ;
        RECT 41.730 51.885 42.020 53.945 ;
        RECT 44.515 52.485 44.990 55.535 ;
        RECT 49.470 52.395 49.880 55.490 ;
        RECT 48.510 50.735 48.820 50.765 ;
        RECT 41.650 44.030 41.975 46.400 ;
        RECT 43.300 46.075 43.700 50.040 ;
        RECT 42.385 40.290 42.730 42.750 ;
        RECT 44.020 41.970 44.345 44.735 ;
        RECT 45.005 44.005 45.410 47.335 ;
        RECT 48.510 44.635 48.825 50.735 ;
        RECT 49.655 41.030 50.025 50.130 ;
        RECT 50.600 42.095 50.890 53.930 ;
        RECT 54.050 52.370 54.460 55.465 ;
        RECT 58.505 51.825 58.815 54.340 ;
        RECT 51.495 44.590 51.825 50.785 ;
        RECT 54.415 44.060 54.855 47.335 ;
        RECT 56.795 46.075 57.320 50.015 ;
        RECT 55.955 41.970 56.280 44.735 ;
        RECT 58.470 44.065 58.885 46.455 ;
        RECT 59.500 42.625 59.815 53.310 ;
        RECT 60.830 47.015 61.315 50.025 ;
        RECT 62.010 42.640 62.340 53.335 ;
        RECT 60.200 41.235 60.535 42.585 ;
        RECT -78.220 22.230 -77.905 33.280 ;
        RECT -74.385 32.575 -73.985 35.625 ;
        RECT -69.465 32.485 -69.055 35.580 ;
        RECT -64.885 32.460 -64.475 35.555 ;
        RECT -76.550 20.380 -76.205 22.840 ;
        RECT -59.435 22.715 -59.120 33.400 ;
        RECT -55.745 25.510 -55.330 28.325 ;
        RECT -55.005 27.095 -54.620 28.990 ;
        RECT -0.030 25.235 0.325 39.175 ;
        RECT 63.315 38.545 63.765 48.810 ;
        RECT 1.595 26.025 1.955 37.575 ;
        RECT 64.480 37.005 64.965 45.890 ;
        RECT 71.420 36.280 71.825 48.325 ;
        RECT 73.495 38.180 73.885 49.605 ;
        RECT 76.655 42.020 77.010 53.105 ;
        RECT 80.400 51.745 80.690 53.805 ;
        RECT 83.170 52.345 83.670 55.395 ;
        RECT 88.140 52.255 88.550 55.350 ;
        RECT 87.180 50.595 87.490 50.625 ;
        RECT 77.980 46.875 78.450 49.865 ;
        RECT 80.330 43.890 80.645 46.260 ;
        RECT 81.950 45.935 82.370 49.900 ;
        RECT 78.615 41.180 78.995 42.555 ;
        RECT 81.055 40.150 81.400 42.610 ;
        RECT 82.690 41.830 83.015 44.595 ;
        RECT 83.675 43.865 84.080 47.195 ;
        RECT 87.180 44.495 87.495 50.595 ;
        RECT 88.325 40.890 88.695 49.990 ;
        RECT 89.270 41.955 89.560 53.790 ;
        RECT 92.720 52.230 93.130 55.325 ;
        RECT 97.175 51.685 97.485 54.200 ;
        RECT 101.425 53.385 101.805 53.765 ;
        RECT 103.555 53.385 103.935 53.765 ;
        RECT 90.165 44.450 90.495 50.645 ;
        RECT 93.070 43.920 93.525 47.195 ;
        RECT 95.430 45.935 95.975 49.875 ;
        RECT 99.485 46.875 99.920 49.885 ;
        RECT 94.625 41.830 94.950 44.595 ;
        RECT 97.140 43.925 97.555 46.315 ;
        RECT 100.680 42.500 101.010 53.195 ;
        RECT 102.115 46.835 102.500 52.620 ;
        RECT 98.870 41.095 99.205 42.445 ;
        RECT 102.475 42.080 102.900 46.355 ;
        RECT 104.175 43.845 104.475 50.885 ;
        RECT 105.295 43.240 105.595 50.170 ;
        RECT 106.605 43.840 106.905 50.190 ;
        RECT 101.135 41.170 101.515 41.550 ;
        RECT 103.330 41.155 103.710 41.535 ;
        RECT 107.200 41.095 107.490 50.875 ;
        RECT 107.920 43.870 108.215 50.695 ;
        RECT 109.050 43.330 109.350 50.140 ;
        RECT 109.840 43.925 110.150 53.965 ;
        RECT 119.030 52.210 119.410 52.590 ;
        RECT 110.635 43.855 110.935 50.685 ;
        RECT 111.760 43.240 112.060 50.180 ;
        RECT 113.210 43.115 113.490 46.150 ;
        RECT 113.970 43.815 114.250 50.175 ;
        RECT 114.820 43.815 115.120 50.635 ;
        RECT 115.960 43.070 116.260 50.225 ;
        RECT 116.605 47.260 116.985 47.640 ;
        RECT 116.605 45.205 116.985 45.585 ;
        RECT 118.455 45.085 118.770 49.410 ;
        RECT 119.065 47.160 119.345 48.690 ;
        RECT 119.635 43.845 119.935 50.885 ;
        RECT 120.755 43.240 121.055 50.170 ;
        RECT 121.410 44.600 121.710 48.660 ;
        RECT 122.065 43.840 122.365 50.190 ;
        RECT 118.930 42.035 119.310 42.415 ;
        RECT 122.660 41.630 122.950 50.875 ;
        RECT 123.380 43.870 123.675 50.695 ;
        RECT 124.510 43.330 124.810 50.140 ;
        RECT 125.300 43.925 125.610 52.660 ;
        RECT 126.095 43.855 126.395 50.685 ;
        RECT 127.220 43.240 127.520 50.180 ;
        RECT 127.900 44.585 128.180 48.675 ;
        RECT 128.670 43.115 128.950 46.150 ;
        RECT 129.430 43.815 129.710 50.175 ;
        RECT 130.280 43.815 130.580 50.635 ;
        RECT 131.420 43.070 131.720 50.225 ;
        RECT 133.760 48.840 134.135 57.040 ;
        RECT 135.505 48.035 135.805 59.030 ;
        RECT 136.490 47.095 136.870 57.350 ;
        RECT 137.360 44.940 137.795 58.515 ;
        RECT 193.070 57.675 193.585 67.975 ;
        RECT 194.755 56.570 195.340 67.350 ;
        RECT 196.240 64.840 196.595 78.760 ;
        RECT 259.585 78.130 260.035 88.395 ;
        RECT 197.865 65.745 198.225 77.160 ;
        RECT 260.750 76.590 261.235 85.475 ;
        RECT 267.415 76.325 267.820 87.855 ;
        RECT 269.490 78.225 269.880 89.325 ;
        RECT 272.915 81.705 273.270 92.790 ;
        RECT 276.660 91.430 276.950 93.490 ;
        RECT 279.430 92.030 279.930 95.080 ;
        RECT 284.400 91.940 284.810 95.035 ;
        RECT 283.440 90.280 283.750 90.310 ;
        RECT 274.240 86.560 274.710 89.550 ;
        RECT 276.590 83.575 276.905 85.945 ;
        RECT 278.210 85.620 278.630 89.585 ;
        RECT 274.875 80.865 275.255 82.240 ;
        RECT 277.315 79.835 277.660 82.295 ;
        RECT 278.950 81.515 279.275 84.280 ;
        RECT 279.935 83.550 280.340 86.880 ;
        RECT 283.440 84.180 283.755 90.280 ;
        RECT 284.585 80.575 284.955 89.675 ;
        RECT 285.530 81.640 285.820 93.475 ;
        RECT 288.980 91.915 289.390 95.010 ;
        RECT 293.435 91.370 293.745 93.885 ;
        RECT 297.685 93.070 298.065 93.450 ;
        RECT 299.815 93.070 300.195 93.450 ;
        RECT 286.425 84.135 286.755 90.330 ;
        RECT 289.330 83.605 289.785 86.880 ;
        RECT 291.690 85.620 292.235 89.560 ;
        RECT 295.745 86.560 296.180 89.570 ;
        RECT 290.885 81.515 291.210 84.280 ;
        RECT 293.400 83.610 293.815 86.000 ;
        RECT 296.940 82.185 297.270 92.880 ;
        RECT 298.375 86.520 298.760 92.305 ;
        RECT 295.130 80.780 295.465 82.130 ;
        RECT 298.735 81.765 299.160 86.040 ;
        RECT 300.435 83.530 300.735 90.570 ;
        RECT 301.555 82.925 301.855 89.855 ;
        RECT 302.865 83.525 303.165 89.875 ;
        RECT 297.395 80.855 297.775 81.235 ;
        RECT 299.590 80.840 299.970 81.220 ;
        RECT 303.460 80.780 303.750 90.560 ;
        RECT 304.180 83.555 304.475 90.380 ;
        RECT 305.310 83.015 305.610 89.825 ;
        RECT 306.100 83.610 306.410 93.650 ;
        RECT 315.290 91.895 315.670 92.275 ;
        RECT 306.895 83.540 307.195 90.370 ;
        RECT 308.020 82.925 308.320 89.865 ;
        RECT 309.470 82.800 309.750 85.835 ;
        RECT 310.230 83.500 310.510 89.860 ;
        RECT 311.080 83.500 311.380 90.320 ;
        RECT 312.220 82.755 312.520 89.910 ;
        RECT 312.865 86.945 313.245 87.325 ;
        RECT 312.865 84.890 313.245 85.270 ;
        RECT 314.715 84.770 315.030 89.095 ;
        RECT 315.325 86.845 315.605 88.375 ;
        RECT 315.895 83.530 316.195 90.570 ;
        RECT 317.015 82.925 317.315 89.855 ;
        RECT 317.670 84.285 317.970 88.345 ;
        RECT 318.325 83.525 318.625 89.875 ;
        RECT 315.190 81.720 315.570 82.100 ;
        RECT 318.920 81.315 319.210 90.560 ;
        RECT 319.640 83.555 319.935 90.380 ;
        RECT 320.770 83.015 321.070 89.825 ;
        RECT 321.560 83.610 321.870 92.345 ;
        RECT 322.355 83.540 322.655 90.370 ;
        RECT 323.480 82.925 323.780 89.865 ;
        RECT 324.160 84.270 324.440 88.360 ;
        RECT 324.930 82.800 325.210 85.835 ;
        RECT 325.690 83.500 325.970 89.860 ;
        RECT 326.540 83.500 326.840 90.320 ;
        RECT 327.680 82.755 327.980 89.910 ;
        RECT 329.965 88.615 330.340 96.900 ;
        RECT 331.710 87.895 332.010 98.890 ;
        RECT 332.880 86.740 333.260 96.995 ;
        RECT 333.750 84.585 334.185 98.160 ;
        RECT 389.455 97.360 389.970 107.410 ;
        RECT 391.140 96.005 391.725 106.785 ;
        RECT 392.990 104.340 393.345 118.130 ;
        RECT 456.335 117.500 456.785 128.000 ;
        RECT 394.615 105.195 394.975 116.530 ;
        RECT 457.500 115.960 457.985 125.200 ;
        RECT 463.915 115.715 464.320 127.245 ;
        RECT 465.990 117.615 466.380 128.715 ;
        RECT 469.395 121.205 469.750 132.290 ;
        RECT 473.140 130.930 473.430 132.990 ;
        RECT 475.910 131.530 476.410 134.580 ;
        RECT 480.880 131.440 481.290 134.535 ;
        RECT 479.920 129.780 480.230 129.810 ;
        RECT 470.720 126.060 471.190 129.050 ;
        RECT 473.070 123.075 473.385 125.445 ;
        RECT 474.690 125.120 475.110 129.085 ;
        RECT 471.355 120.365 471.735 121.740 ;
        RECT 473.795 119.335 474.140 121.795 ;
        RECT 475.430 121.015 475.755 123.780 ;
        RECT 476.415 123.050 476.820 126.380 ;
        RECT 479.920 123.680 480.235 129.780 ;
        RECT 481.065 120.075 481.435 129.175 ;
        RECT 482.010 121.140 482.300 132.975 ;
        RECT 485.460 131.415 485.870 134.510 ;
        RECT 489.915 130.870 490.225 133.385 ;
        RECT 494.165 132.570 494.545 132.950 ;
        RECT 496.295 132.570 496.675 132.950 ;
        RECT 482.905 123.635 483.235 129.830 ;
        RECT 485.810 123.105 486.265 126.380 ;
        RECT 488.170 125.120 488.715 129.060 ;
        RECT 492.225 126.060 492.660 129.070 ;
        RECT 487.365 121.015 487.690 123.780 ;
        RECT 489.880 123.110 490.295 125.500 ;
        RECT 493.420 121.685 493.750 132.380 ;
        RECT 494.855 126.020 495.240 131.805 ;
        RECT 491.610 120.280 491.945 121.630 ;
        RECT 495.215 121.265 495.640 125.540 ;
        RECT 496.915 123.030 497.215 130.070 ;
        RECT 498.035 122.425 498.335 129.355 ;
        RECT 499.345 123.025 499.645 129.375 ;
        RECT 493.875 120.355 494.255 120.735 ;
        RECT 496.070 120.340 496.450 120.720 ;
        RECT 499.940 120.280 500.230 130.060 ;
        RECT 500.660 123.055 500.955 129.880 ;
        RECT 501.790 122.515 502.090 129.325 ;
        RECT 502.580 123.110 502.890 133.150 ;
        RECT 511.770 131.395 512.150 131.775 ;
        RECT 503.375 123.040 503.675 129.870 ;
        RECT 504.500 122.425 504.800 129.365 ;
        RECT 505.950 122.300 506.230 125.335 ;
        RECT 506.710 123.000 506.990 129.360 ;
        RECT 507.560 123.000 507.860 129.820 ;
        RECT 508.700 122.255 509.000 129.410 ;
        RECT 509.345 126.445 509.725 126.825 ;
        RECT 509.345 124.390 509.725 124.770 ;
        RECT 511.195 124.270 511.510 128.595 ;
        RECT 511.805 126.345 512.085 127.875 ;
        RECT 512.375 123.030 512.675 130.070 ;
        RECT 513.495 122.425 513.795 129.355 ;
        RECT 514.150 123.785 514.450 127.845 ;
        RECT 514.805 123.025 515.105 129.375 ;
        RECT 511.670 121.220 512.050 121.600 ;
        RECT 515.400 120.815 515.690 130.060 ;
        RECT 516.120 123.055 516.415 129.880 ;
        RECT 517.250 122.515 517.550 129.325 ;
        RECT 518.040 123.110 518.350 131.845 ;
        RECT 518.835 123.040 519.135 129.870 ;
        RECT 519.960 122.425 520.260 129.365 ;
        RECT 520.640 123.770 520.920 127.860 ;
        RECT 521.410 122.300 521.690 125.335 ;
        RECT 522.170 123.000 522.450 129.360 ;
        RECT 523.020 123.000 523.320 129.820 ;
        RECT 524.160 122.255 524.460 129.410 ;
        RECT 526.345 128.045 526.720 136.245 ;
        RECT 528.090 127.240 528.390 138.235 ;
        RECT 529.200 126.335 529.580 136.590 ;
        RECT 530.070 124.180 530.505 137.755 ;
        RECT 585.775 136.955 586.290 147.005 ;
        RECT 587.460 135.600 588.045 146.380 ;
        RECT 589.155 143.915 589.510 157.705 ;
        RECT 652.500 157.075 652.950 167.340 ;
        RECT 590.780 144.770 591.140 156.105 ;
        RECT 653.665 155.535 654.150 164.420 ;
        RECT 659.970 155.160 660.375 166.690 ;
        RECT 662.045 157.060 662.435 168.160 ;
        RECT 665.815 160.610 666.170 171.695 ;
        RECT 669.560 170.335 669.850 172.395 ;
        RECT 672.330 170.935 672.830 173.985 ;
        RECT 677.300 170.845 677.710 173.940 ;
        RECT 676.340 169.185 676.650 169.215 ;
        RECT 667.140 165.465 667.610 168.455 ;
        RECT 669.490 162.480 669.805 164.850 ;
        RECT 671.110 164.525 671.530 168.490 ;
        RECT 667.775 159.770 668.155 161.145 ;
        RECT 670.215 158.740 670.560 161.200 ;
        RECT 671.850 160.420 672.175 163.185 ;
        RECT 672.835 162.455 673.240 165.785 ;
        RECT 676.340 163.085 676.655 169.185 ;
        RECT 677.485 159.480 677.855 168.580 ;
        RECT 678.430 160.545 678.720 172.380 ;
        RECT 681.880 170.820 682.290 173.915 ;
        RECT 686.335 170.275 686.645 172.790 ;
        RECT 690.585 171.975 690.965 172.355 ;
        RECT 692.715 171.975 693.095 172.355 ;
        RECT 679.325 163.040 679.655 169.235 ;
        RECT 682.230 162.510 682.685 165.785 ;
        RECT 684.590 164.525 685.135 168.465 ;
        RECT 688.645 165.465 689.080 168.475 ;
        RECT 683.785 160.420 684.110 163.185 ;
        RECT 686.300 162.515 686.715 164.905 ;
        RECT 689.840 161.090 690.170 171.785 ;
        RECT 691.275 165.425 691.660 171.210 ;
        RECT 688.030 159.685 688.365 161.035 ;
        RECT 691.635 160.670 692.060 164.945 ;
        RECT 693.335 162.435 693.635 169.475 ;
        RECT 694.455 161.830 694.755 168.760 ;
        RECT 695.765 162.430 696.065 168.780 ;
        RECT 690.295 159.760 690.675 160.140 ;
        RECT 692.490 159.745 692.870 160.125 ;
        RECT 696.360 159.685 696.650 169.465 ;
        RECT 697.080 162.460 697.375 169.285 ;
        RECT 698.210 161.920 698.510 168.730 ;
        RECT 699.000 162.515 699.310 172.555 ;
        RECT 708.190 170.800 708.570 171.180 ;
        RECT 699.795 162.445 700.095 169.275 ;
        RECT 700.920 161.830 701.220 168.770 ;
        RECT 702.370 161.705 702.650 164.740 ;
        RECT 703.130 162.405 703.410 168.765 ;
        RECT 703.980 162.405 704.280 169.225 ;
        RECT 705.120 161.660 705.420 168.815 ;
        RECT 705.765 165.850 706.145 166.230 ;
        RECT 705.765 163.795 706.145 164.175 ;
        RECT 707.615 163.675 707.930 168.000 ;
        RECT 708.225 165.750 708.505 167.280 ;
        RECT 708.795 162.435 709.095 169.475 ;
        RECT 710.570 163.190 710.870 167.250 ;
        RECT 708.090 160.625 708.470 161.005 ;
        RECT 711.820 160.220 712.110 169.465 ;
        RECT 713.670 161.920 713.970 168.730 ;
        RECT 714.460 162.515 714.770 171.250 ;
        RECT 715.255 162.445 715.555 169.275 ;
        RECT 717.060 163.175 717.340 167.265 ;
        RECT 717.830 161.705 718.110 164.740 ;
        RECT 720.580 161.660 720.880 168.815 ;
        RECT 757.410 160.705 757.725 171.755 ;
        RECT 761.245 171.050 761.645 174.100 ;
        RECT 766.165 170.960 766.575 174.055 ;
        RECT 770.745 170.935 771.155 174.030 ;
        RECT 759.080 158.855 759.425 161.315 ;
        RECT 776.195 161.190 776.510 171.875 ;
        RECT 781.380 163.980 781.830 168.140 ;
        RECT 790.815 167.670 791.195 168.050 ;
        RECT 783.080 166.960 783.605 167.400 ;
        RECT 790.805 166.920 791.185 167.300 ;
        RECT 594.430 147.980 594.810 148.360 ;
        RECT 594.420 147.230 594.800 147.610 ;
        RECT 594.465 146.545 594.845 146.925 ;
        RECT 594.430 145.875 594.810 146.255 ;
        RECT 595.145 142.800 595.445 149.840 ;
        RECT 596.265 142.195 596.565 149.125 ;
        RECT 596.920 143.555 597.220 147.615 ;
        RECT 597.575 142.795 597.875 149.145 ;
        RECT 598.170 144.670 598.490 149.830 ;
        RECT 598.890 142.825 599.185 149.650 ;
        RECT 600.020 142.285 600.320 149.095 ;
        RECT 600.810 142.880 601.120 149.070 ;
        RECT 601.605 142.810 601.905 149.640 ;
        RECT 602.730 142.195 603.030 149.135 ;
        RECT 603.410 143.540 603.690 147.630 ;
        RECT 604.180 142.070 604.460 145.105 ;
        RECT 604.940 142.770 605.245 149.130 ;
        RECT 605.790 142.770 606.090 149.590 ;
        RECT 606.930 142.025 607.230 149.180 ;
        RECT 607.595 147.980 607.975 148.360 ;
        RECT 609.865 147.980 610.245 148.385 ;
        RECT 607.600 147.230 607.980 147.610 ;
        RECT 609.870 147.230 610.250 147.635 ;
        RECT 607.600 146.215 607.980 146.595 ;
        RECT 609.385 144.795 609.705 146.925 ;
        RECT 607.815 141.505 608.195 144.525 ;
        RECT 609.995 143.955 610.275 146.360 ;
        RECT 610.605 142.800 610.905 149.840 ;
        RECT 611.725 142.195 612.025 149.125 ;
        RECT 612.380 143.555 612.680 147.615 ;
        RECT 613.035 142.795 613.335 149.145 ;
        RECT 613.630 144.670 613.955 149.830 ;
        RECT 614.350 142.825 614.645 149.650 ;
        RECT 615.480 142.285 615.780 149.095 ;
        RECT 616.270 142.880 616.580 149.070 ;
        RECT 617.065 142.810 617.365 149.640 ;
        RECT 618.190 142.195 618.490 149.135 ;
        RECT 618.870 143.540 619.150 147.630 ;
        RECT 619.640 142.070 619.920 145.105 ;
        RECT 620.400 142.770 620.720 149.130 ;
        RECT 621.250 142.770 621.550 149.590 ;
        RECT 622.390 142.025 622.690 149.180 ;
        RECT 623.330 147.980 623.690 149.810 ;
        RECT 623.025 144.170 623.405 144.550 ;
        RECT 623.730 140.055 624.090 146.615 ;
        RECT 624.870 144.805 625.195 146.670 ;
        RECT 625.510 146.460 625.925 149.810 ;
        RECT 625.535 141.460 625.995 146.145 ;
        RECT 626.320 144.005 626.770 152.825 ;
        RECT 627.180 141.630 627.535 151.935 ;
        RECT 627.845 147.235 628.190 148.290 ;
        RECT 628.505 145.830 628.935 148.820 ;
        RECT 626.250 140.115 626.630 140.495 ;
        RECT 629.140 140.135 629.520 141.510 ;
        RECT 629.910 140.955 630.225 152.005 ;
        RECT 630.925 150.700 631.215 152.760 ;
        RECT 633.710 151.300 634.185 154.350 ;
        RECT 638.665 151.210 639.075 154.305 ;
        RECT 637.705 149.550 638.015 149.580 ;
        RECT 630.845 142.845 631.170 145.215 ;
        RECT 632.495 144.890 632.895 148.855 ;
        RECT 631.580 139.105 631.925 141.565 ;
        RECT 633.215 140.785 633.540 143.550 ;
        RECT 634.200 142.820 634.605 146.150 ;
        RECT 637.705 143.450 638.020 149.550 ;
        RECT 638.850 139.845 639.220 148.945 ;
        RECT 639.795 140.910 640.085 152.745 ;
        RECT 643.245 151.185 643.655 154.280 ;
        RECT 647.700 150.640 648.010 153.155 ;
        RECT 640.690 143.405 641.020 149.600 ;
        RECT 643.610 142.875 644.050 146.150 ;
        RECT 645.990 144.890 646.515 148.830 ;
        RECT 645.150 140.785 645.475 143.550 ;
        RECT 647.665 142.880 648.080 145.270 ;
        RECT 648.695 141.440 649.010 152.125 ;
        RECT 650.025 145.830 650.510 148.840 ;
        RECT 651.205 141.455 651.535 152.150 ;
        RECT 649.395 140.050 649.730 141.400 ;
        RECT 561.020 121.180 561.335 132.230 ;
        RECT 564.855 131.525 565.255 134.575 ;
        RECT 569.775 131.435 570.185 134.530 ;
        RECT 574.355 131.410 574.765 134.505 ;
        RECT 562.690 119.330 563.035 121.790 ;
        RECT 579.805 121.665 580.120 132.350 ;
        RECT 584.990 124.455 585.440 128.615 ;
        RECT 586.690 127.435 587.215 127.875 ;
        RECT 398.050 108.395 398.430 108.775 ;
        RECT 398.040 107.645 398.420 108.025 ;
        RECT 398.085 106.960 398.465 107.340 ;
        RECT 398.050 106.290 398.430 106.670 ;
        RECT 398.765 103.215 399.065 110.255 ;
        RECT 399.885 102.610 400.185 109.540 ;
        RECT 400.540 103.970 400.840 108.030 ;
        RECT 401.195 103.210 401.495 109.560 ;
        RECT 401.790 105.085 402.110 110.245 ;
        RECT 402.510 103.240 402.805 110.065 ;
        RECT 403.640 102.700 403.940 109.510 ;
        RECT 404.430 103.295 404.740 109.485 ;
        RECT 405.225 103.225 405.525 110.055 ;
        RECT 406.350 102.610 406.650 109.550 ;
        RECT 407.030 103.955 407.310 108.045 ;
        RECT 407.800 102.485 408.080 105.520 ;
        RECT 408.560 103.185 408.865 109.545 ;
        RECT 409.410 103.185 409.710 110.005 ;
        RECT 410.550 102.440 410.850 109.595 ;
        RECT 411.215 108.395 411.595 108.775 ;
        RECT 413.485 108.395 413.865 108.800 ;
        RECT 411.220 107.645 411.600 108.025 ;
        RECT 413.490 107.645 413.870 108.050 ;
        RECT 411.220 106.630 411.600 107.010 ;
        RECT 413.005 105.210 413.325 107.340 ;
        RECT 411.435 101.920 411.815 104.940 ;
        RECT 413.615 104.370 413.895 106.775 ;
        RECT 414.225 103.215 414.525 110.255 ;
        RECT 415.345 102.610 415.645 109.540 ;
        RECT 416.000 103.970 416.300 108.030 ;
        RECT 416.655 103.210 416.955 109.560 ;
        RECT 417.250 105.085 417.575 110.245 ;
        RECT 417.970 103.240 418.265 110.065 ;
        RECT 419.100 102.700 419.400 109.510 ;
        RECT 419.890 103.295 420.200 109.485 ;
        RECT 420.685 103.225 420.985 110.055 ;
        RECT 421.810 102.610 422.110 109.550 ;
        RECT 422.490 103.955 422.770 108.045 ;
        RECT 423.260 102.485 423.540 105.520 ;
        RECT 424.020 103.185 424.340 109.545 ;
        RECT 424.870 103.185 425.170 110.005 ;
        RECT 426.010 102.440 426.310 109.595 ;
        RECT 426.950 108.395 427.310 110.225 ;
        RECT 426.645 104.585 427.025 104.965 ;
        RECT 427.350 100.470 427.710 107.030 ;
        RECT 428.490 105.220 428.815 107.085 ;
        RECT 429.130 106.875 429.545 110.225 ;
        RECT 429.155 101.875 429.615 106.560 ;
        RECT 429.940 104.420 430.390 113.240 ;
        RECT 430.800 102.045 431.155 112.350 ;
        RECT 431.465 107.650 431.810 108.705 ;
        RECT 432.125 106.245 432.555 109.235 ;
        RECT 429.870 100.530 430.250 100.910 ;
        RECT 432.760 100.550 433.140 101.925 ;
        RECT 433.530 101.370 433.845 112.420 ;
        RECT 434.545 111.115 434.835 113.175 ;
        RECT 437.330 111.715 437.805 114.765 ;
        RECT 442.285 111.625 442.695 114.720 ;
        RECT 441.325 109.965 441.635 109.995 ;
        RECT 434.465 103.260 434.790 105.630 ;
        RECT 436.115 105.305 436.515 109.270 ;
        RECT 435.200 99.520 435.545 101.980 ;
        RECT 436.835 101.200 437.160 103.965 ;
        RECT 437.820 103.235 438.225 106.565 ;
        RECT 441.325 103.865 441.640 109.965 ;
        RECT 442.470 100.260 442.840 109.360 ;
        RECT 443.415 101.325 443.705 113.160 ;
        RECT 446.865 111.600 447.275 114.695 ;
        RECT 451.320 111.055 451.630 113.570 ;
        RECT 444.310 103.820 444.640 110.015 ;
        RECT 447.230 103.290 447.670 106.565 ;
        RECT 449.610 105.305 450.135 109.245 ;
        RECT 448.770 101.200 449.095 103.965 ;
        RECT 451.285 103.295 451.700 105.685 ;
        RECT 452.315 101.855 452.630 112.540 ;
        RECT 453.645 106.245 454.130 109.255 ;
        RECT 454.825 101.870 455.155 112.565 ;
        RECT 453.015 100.465 453.350 101.815 ;
        RECT 364.660 81.640 364.975 92.690 ;
        RECT 368.495 91.985 368.895 95.035 ;
        RECT 373.415 91.895 373.825 94.990 ;
        RECT 377.995 91.870 378.405 94.965 ;
        RECT 366.330 79.790 366.675 82.250 ;
        RECT 383.445 82.125 383.760 92.810 ;
        RECT 388.630 84.915 389.080 89.075 ;
        RECT 390.330 87.895 390.855 88.335 ;
        RECT 201.650 68.975 202.030 69.355 ;
        RECT 201.640 68.225 202.020 68.605 ;
        RECT 201.685 67.540 202.065 67.920 ;
        RECT 201.650 66.870 202.030 67.250 ;
        RECT 202.365 63.795 202.665 70.835 ;
        RECT 203.485 63.190 203.785 70.120 ;
        RECT 204.140 64.550 204.440 68.610 ;
        RECT 204.795 63.790 205.095 70.140 ;
        RECT 205.390 65.665 205.710 70.825 ;
        RECT 206.110 63.820 206.405 70.645 ;
        RECT 207.240 63.280 207.540 70.090 ;
        RECT 208.030 63.875 208.340 70.065 ;
        RECT 208.825 63.805 209.125 70.635 ;
        RECT 209.950 63.190 210.250 70.130 ;
        RECT 210.630 64.535 210.910 68.625 ;
        RECT 211.400 63.065 211.680 66.100 ;
        RECT 212.160 63.765 212.465 70.125 ;
        RECT 213.010 63.765 213.310 70.585 ;
        RECT 214.150 63.020 214.450 70.175 ;
        RECT 214.815 68.975 215.195 69.355 ;
        RECT 217.085 68.975 217.465 69.380 ;
        RECT 214.820 68.225 215.200 68.605 ;
        RECT 217.090 68.225 217.470 68.630 ;
        RECT 214.820 67.210 215.200 67.590 ;
        RECT 216.605 65.790 216.925 67.920 ;
        RECT 215.035 62.500 215.415 65.520 ;
        RECT 217.215 64.950 217.495 67.355 ;
        RECT 217.825 63.795 218.125 70.835 ;
        RECT 218.945 63.190 219.245 70.120 ;
        RECT 219.600 64.550 219.900 68.610 ;
        RECT 220.255 63.790 220.555 70.140 ;
        RECT 220.850 65.665 221.175 70.825 ;
        RECT 221.570 63.820 221.865 70.645 ;
        RECT 222.700 63.280 223.000 70.090 ;
        RECT 223.490 63.875 223.800 70.065 ;
        RECT 224.285 63.805 224.585 70.635 ;
        RECT 225.410 63.190 225.710 70.130 ;
        RECT 226.090 64.535 226.370 68.625 ;
        RECT 226.860 63.065 227.140 66.100 ;
        RECT 227.620 63.765 227.940 70.125 ;
        RECT 228.470 63.765 228.770 70.585 ;
        RECT 229.610 63.020 229.910 70.175 ;
        RECT 230.550 68.975 230.910 70.805 ;
        RECT 230.245 65.165 230.625 65.545 ;
        RECT 230.950 61.050 231.310 67.610 ;
        RECT 232.090 65.800 232.415 67.665 ;
        RECT 232.730 67.455 233.145 70.805 ;
        RECT 232.755 62.455 233.215 67.140 ;
        RECT 233.540 65.000 233.990 73.820 ;
        RECT 234.400 62.625 234.755 72.930 ;
        RECT 235.065 68.230 235.410 69.285 ;
        RECT 235.725 66.825 236.155 69.815 ;
        RECT 233.470 61.110 233.850 61.490 ;
        RECT 236.360 61.130 236.740 62.505 ;
        RECT 237.130 61.950 237.445 73.000 ;
        RECT 238.145 71.695 238.435 73.755 ;
        RECT 240.930 72.295 241.405 75.345 ;
        RECT 245.885 72.205 246.295 75.300 ;
        RECT 244.925 70.545 245.235 70.575 ;
        RECT 238.065 63.840 238.390 66.210 ;
        RECT 239.715 65.885 240.115 69.850 ;
        RECT 238.800 60.100 239.145 62.560 ;
        RECT 240.435 61.780 240.760 64.545 ;
        RECT 241.420 63.815 241.825 67.145 ;
        RECT 244.925 64.445 245.240 70.545 ;
        RECT 246.070 60.840 246.440 69.940 ;
        RECT 247.015 61.905 247.305 73.740 ;
        RECT 250.465 72.180 250.875 75.275 ;
        RECT 254.920 71.635 255.230 74.150 ;
        RECT 247.910 64.400 248.240 70.595 ;
        RECT 250.830 63.870 251.270 67.145 ;
        RECT 253.210 65.885 253.735 69.825 ;
        RECT 252.370 61.780 252.695 64.545 ;
        RECT 254.885 63.875 255.300 66.265 ;
        RECT 255.915 62.435 256.230 73.120 ;
        RECT 257.245 66.825 257.730 69.835 ;
        RECT 258.425 62.450 258.755 73.145 ;
        RECT 256.615 61.045 256.950 62.395 ;
        RECT 168.270 42.130 168.585 53.180 ;
        RECT 172.105 52.475 172.505 55.525 ;
        RECT 177.025 52.385 177.435 55.480 ;
        RECT 181.605 52.360 182.015 55.455 ;
        RECT 169.940 40.280 170.285 42.740 ;
        RECT 187.055 42.615 187.370 53.300 ;
        RECT 192.240 45.405 192.690 49.565 ;
        RECT 193.940 48.385 194.465 48.825 ;
        RECT 5.240 27.935 5.620 28.315 ;
        RECT 5.205 27.265 5.585 27.645 ;
        RECT 5.920 24.190 6.220 31.230 ;
        RECT 7.040 23.585 7.340 30.515 ;
        RECT 8.350 24.185 8.650 30.535 ;
        RECT 8.945 26.060 9.265 31.220 ;
        RECT 9.665 24.215 9.960 31.040 ;
        RECT 10.795 23.675 11.095 30.485 ;
        RECT 11.585 24.270 11.895 30.460 ;
        RECT 12.380 24.200 12.680 31.030 ;
        RECT 13.505 23.585 13.805 30.525 ;
        RECT 14.955 23.460 15.235 26.495 ;
        RECT 15.715 24.160 16.020 30.520 ;
        RECT 16.565 24.160 16.865 30.980 ;
        RECT 17.705 23.415 18.005 30.570 ;
        RECT 18.375 27.605 18.755 27.985 ;
        RECT 20.160 26.185 20.480 28.315 ;
        RECT 18.590 22.895 18.970 25.915 ;
        RECT 20.770 25.345 21.050 27.750 ;
        RECT 21.380 24.190 21.680 31.230 ;
        RECT 22.500 23.585 22.800 30.515 ;
        RECT 23.810 24.185 24.110 30.535 ;
        RECT 24.405 26.060 24.730 31.220 ;
        RECT 25.125 24.215 25.420 31.040 ;
        RECT 26.255 23.675 26.555 30.485 ;
        RECT 27.045 24.270 27.355 30.460 ;
        RECT 27.840 24.200 28.140 31.030 ;
        RECT 28.965 23.585 29.265 30.525 ;
        RECT 30.415 23.460 30.695 26.495 ;
        RECT 31.175 24.160 31.495 30.520 ;
        RECT 32.025 24.160 32.325 30.980 ;
        RECT 33.165 23.415 33.465 30.570 ;
        RECT 33.800 25.560 34.180 25.940 ;
        RECT 34.505 21.445 34.865 28.005 ;
        RECT 35.645 26.195 35.970 28.060 ;
        RECT 36.310 22.850 36.770 27.535 ;
        RECT 37.095 25.395 37.545 34.215 ;
        RECT 39.280 27.220 39.710 30.210 ;
        RECT 37.025 21.505 37.405 21.885 ;
        RECT 39.915 21.525 40.295 22.900 ;
        RECT 40.685 22.345 41.000 33.395 ;
        RECT 41.700 32.090 41.990 34.150 ;
        RECT 44.485 32.690 44.960 35.740 ;
        RECT 49.440 32.600 49.850 35.695 ;
        RECT 41.620 24.235 41.945 26.605 ;
        RECT 43.270 26.280 43.670 30.245 ;
        RECT 42.355 20.495 42.700 22.955 ;
        RECT 43.990 22.175 44.315 24.940 ;
        RECT 44.975 24.210 45.380 27.540 ;
        RECT 49.625 21.235 49.995 30.335 ;
        RECT 50.570 22.300 50.860 34.135 ;
        RECT 54.020 32.575 54.430 35.670 ;
        RECT 58.475 32.030 58.785 34.545 ;
        RECT 54.385 24.265 54.825 27.540 ;
        RECT 56.765 26.280 57.290 30.220 ;
        RECT 55.925 22.175 56.250 24.940 ;
        RECT 58.440 24.270 58.855 26.660 ;
        RECT 59.470 22.830 59.785 33.515 ;
        RECT 60.800 27.220 61.285 30.230 ;
        RECT 67.260 29.140 70.585 29.730 ;
        RECT 67.260 28.525 68.010 29.140 ;
        RECT 69.165 25.685 69.835 28.335 ;
        RECT 60.170 21.440 60.505 22.790 ;
        RECT 71.125 9.530 71.575 28.570 ;
        RECT 72.915 8.755 73.330 29.935 ;
        RECT 76.655 22.355 77.010 33.440 ;
        RECT 80.400 32.080 80.690 34.140 ;
        RECT 83.170 32.680 83.670 35.730 ;
        RECT 88.140 32.590 88.550 35.685 ;
        RECT 87.180 30.930 87.490 30.960 ;
        RECT 77.980 27.210 78.450 30.200 ;
        RECT 80.330 24.225 80.645 26.595 ;
        RECT 81.950 26.270 82.370 30.235 ;
        RECT 78.615 21.515 78.995 22.890 ;
        RECT 81.055 20.485 81.400 22.945 ;
        RECT 82.690 22.165 83.015 24.930 ;
        RECT 83.675 24.200 84.080 27.530 ;
        RECT 87.180 24.830 87.495 30.930 ;
        RECT 88.325 21.225 88.695 30.325 ;
        RECT 89.270 22.290 89.560 34.125 ;
        RECT 92.720 32.565 93.130 35.660 ;
        RECT 97.175 32.020 97.485 34.535 ;
        RECT 101.425 33.720 101.805 34.100 ;
        RECT 103.555 33.720 103.935 34.100 ;
        RECT 90.165 24.785 90.495 30.980 ;
        RECT 93.070 24.255 93.525 27.530 ;
        RECT 95.430 26.270 95.975 30.210 ;
        RECT 99.485 27.210 99.920 30.220 ;
        RECT 94.625 22.165 94.950 24.930 ;
        RECT 97.140 24.260 97.555 26.650 ;
        RECT 100.680 22.835 101.010 33.530 ;
        RECT 102.115 27.170 102.500 32.955 ;
        RECT 98.870 21.430 99.205 22.780 ;
        RECT 102.475 22.415 102.900 26.690 ;
        RECT 104.175 24.180 104.475 31.220 ;
        RECT 105.295 23.575 105.595 30.505 ;
        RECT 106.605 24.175 106.905 30.525 ;
        RECT 101.135 21.505 101.515 21.885 ;
        RECT 103.330 21.490 103.710 21.870 ;
        RECT 107.200 21.430 107.490 31.210 ;
        RECT 107.920 24.205 108.215 31.030 ;
        RECT 109.050 23.665 109.350 30.475 ;
        RECT 109.840 24.260 110.150 34.300 ;
        RECT 119.030 32.545 119.410 32.925 ;
        RECT 110.635 24.190 110.935 31.020 ;
        RECT 111.760 23.575 112.060 30.515 ;
        RECT 113.210 23.450 113.490 26.485 ;
        RECT 113.970 24.150 114.250 30.510 ;
        RECT 114.820 24.150 115.120 30.970 ;
        RECT 115.960 23.405 116.260 30.560 ;
        RECT 116.605 27.595 116.985 27.975 ;
        RECT 116.605 25.540 116.985 25.920 ;
        RECT 118.455 25.420 118.770 29.745 ;
        RECT 119.065 27.495 119.345 29.025 ;
        RECT 119.635 24.180 119.935 31.220 ;
        RECT 120.755 23.575 121.055 30.505 ;
        RECT 121.410 24.935 121.710 28.995 ;
        RECT 122.065 24.175 122.365 30.525 ;
        RECT 118.930 22.370 119.310 22.750 ;
        RECT 122.660 21.965 122.950 31.210 ;
        RECT 123.380 24.205 123.675 31.030 ;
        RECT 124.510 23.665 124.810 30.475 ;
        RECT 125.300 24.260 125.610 32.995 ;
        RECT 126.095 24.190 126.395 31.020 ;
        RECT 127.220 23.575 127.520 30.515 ;
        RECT 127.900 24.920 128.180 29.010 ;
        RECT 128.670 23.450 128.950 26.485 ;
        RECT 129.430 24.150 129.710 30.510 ;
        RECT 130.280 24.150 130.580 30.970 ;
        RECT 131.420 23.405 131.720 30.560 ;
        RECT 133.345 29.325 133.720 37.165 ;
        RECT 135.200 28.575 135.500 39.115 ;
        RECT 136.490 27.435 136.870 37.690 ;
        RECT 137.360 25.280 137.795 38.855 ;
        RECT 193.070 38.120 193.585 48.170 ;
        RECT 194.755 36.765 195.340 47.545 ;
        RECT 196.335 45.075 196.690 58.985 ;
        RECT 259.680 58.355 260.130 68.620 ;
        RECT 197.960 45.995 198.320 57.385 ;
        RECT 260.845 56.815 261.330 65.700 ;
        RECT 267.675 56.170 268.080 68.050 ;
        RECT 269.750 58.070 270.140 69.650 ;
        RECT 273.020 61.990 273.375 73.075 ;
        RECT 276.765 71.715 277.055 73.775 ;
        RECT 279.535 72.315 280.035 75.365 ;
        RECT 284.505 72.225 284.915 75.320 ;
        RECT 283.545 70.565 283.855 70.595 ;
        RECT 274.345 66.845 274.815 69.835 ;
        RECT 276.695 63.860 277.010 66.230 ;
        RECT 278.315 65.905 278.735 69.870 ;
        RECT 274.980 61.150 275.360 62.525 ;
        RECT 277.420 60.120 277.765 62.580 ;
        RECT 279.055 61.800 279.380 64.565 ;
        RECT 280.040 63.835 280.445 67.165 ;
        RECT 283.545 64.465 283.860 70.565 ;
        RECT 284.690 60.860 285.060 69.960 ;
        RECT 285.635 61.925 285.925 73.760 ;
        RECT 289.085 72.200 289.495 75.295 ;
        RECT 293.540 71.655 293.850 74.170 ;
        RECT 297.790 73.355 298.170 73.735 ;
        RECT 299.920 73.355 300.300 73.735 ;
        RECT 286.530 64.420 286.860 70.615 ;
        RECT 289.435 63.890 289.890 67.165 ;
        RECT 291.795 65.905 292.340 69.845 ;
        RECT 295.850 66.845 296.285 69.855 ;
        RECT 290.990 61.800 291.315 64.565 ;
        RECT 293.505 63.895 293.920 66.285 ;
        RECT 297.045 62.470 297.375 73.165 ;
        RECT 298.480 66.805 298.865 72.590 ;
        RECT 295.235 61.065 295.570 62.415 ;
        RECT 298.840 62.050 299.265 66.325 ;
        RECT 300.540 63.815 300.840 70.855 ;
        RECT 301.660 63.210 301.960 70.140 ;
        RECT 302.970 63.810 303.270 70.160 ;
        RECT 297.500 61.140 297.880 61.520 ;
        RECT 299.695 61.125 300.075 61.505 ;
        RECT 303.565 61.065 303.855 70.845 ;
        RECT 304.285 63.840 304.580 70.665 ;
        RECT 305.415 63.300 305.715 70.110 ;
        RECT 306.205 63.895 306.515 73.935 ;
        RECT 315.395 72.180 315.775 72.560 ;
        RECT 307.000 63.825 307.300 70.655 ;
        RECT 308.125 63.210 308.425 70.150 ;
        RECT 309.575 63.085 309.855 66.120 ;
        RECT 310.335 63.785 310.615 70.145 ;
        RECT 311.185 63.785 311.485 70.605 ;
        RECT 312.325 63.040 312.625 70.195 ;
        RECT 312.970 67.230 313.350 67.610 ;
        RECT 312.970 65.175 313.350 65.555 ;
        RECT 314.820 65.055 315.135 69.380 ;
        RECT 315.430 67.130 315.710 68.660 ;
        RECT 316.000 63.815 316.300 70.855 ;
        RECT 317.120 63.210 317.420 70.140 ;
        RECT 317.775 64.570 318.075 68.630 ;
        RECT 318.430 63.810 318.730 70.160 ;
        RECT 315.295 62.005 315.675 62.385 ;
        RECT 319.025 61.600 319.315 70.845 ;
        RECT 319.745 63.840 320.040 70.665 ;
        RECT 320.875 63.300 321.175 70.110 ;
        RECT 321.665 63.895 321.975 72.630 ;
        RECT 322.460 63.825 322.760 70.655 ;
        RECT 323.585 63.210 323.885 70.150 ;
        RECT 324.265 64.555 324.545 68.645 ;
        RECT 325.035 63.085 325.315 66.120 ;
        RECT 325.795 63.785 326.075 70.145 ;
        RECT 326.645 63.785 326.945 70.605 ;
        RECT 327.785 63.040 328.085 70.195 ;
        RECT 329.865 68.915 330.240 77.195 ;
        RECT 331.610 68.075 331.910 79.185 ;
        RECT 332.880 67.030 333.260 77.285 ;
        RECT 333.750 64.875 334.185 78.450 ;
        RECT 389.460 77.650 389.975 87.700 ;
        RECT 391.145 76.295 391.730 87.075 ;
        RECT 392.945 84.550 393.300 98.340 ;
        RECT 456.290 97.710 456.740 108.200 ;
        RECT 394.570 85.455 394.930 96.740 ;
        RECT 457.455 96.170 457.940 105.330 ;
        RECT 463.915 95.980 464.320 107.510 ;
        RECT 465.990 97.880 466.380 108.980 ;
        RECT 469.395 101.410 469.750 112.495 ;
        RECT 473.140 111.135 473.430 113.195 ;
        RECT 475.910 111.735 476.410 114.785 ;
        RECT 480.880 111.645 481.290 114.740 ;
        RECT 479.920 109.985 480.230 110.015 ;
        RECT 470.720 106.265 471.190 109.255 ;
        RECT 473.070 103.280 473.385 105.650 ;
        RECT 474.690 105.325 475.110 109.290 ;
        RECT 471.355 100.570 471.735 101.945 ;
        RECT 473.795 99.540 474.140 102.000 ;
        RECT 475.430 101.220 475.755 103.985 ;
        RECT 476.415 103.255 476.820 106.585 ;
        RECT 479.920 103.885 480.235 109.985 ;
        RECT 481.065 100.280 481.435 109.380 ;
        RECT 482.010 101.345 482.300 113.180 ;
        RECT 485.460 111.620 485.870 114.715 ;
        RECT 489.915 111.075 490.225 113.590 ;
        RECT 494.165 112.775 494.545 113.155 ;
        RECT 496.295 112.775 496.675 113.155 ;
        RECT 482.905 103.840 483.235 110.035 ;
        RECT 485.810 103.310 486.265 106.585 ;
        RECT 488.170 105.325 488.715 109.265 ;
        RECT 492.225 106.265 492.660 109.275 ;
        RECT 487.365 101.220 487.690 103.985 ;
        RECT 489.880 103.315 490.295 105.705 ;
        RECT 493.420 101.890 493.750 112.585 ;
        RECT 494.855 106.225 495.240 112.010 ;
        RECT 491.610 100.485 491.945 101.835 ;
        RECT 495.215 101.470 495.640 105.745 ;
        RECT 496.915 103.235 497.215 110.275 ;
        RECT 498.035 102.630 498.335 109.560 ;
        RECT 499.345 103.230 499.645 109.580 ;
        RECT 493.875 100.560 494.255 100.940 ;
        RECT 496.070 100.545 496.450 100.925 ;
        RECT 499.940 100.485 500.230 110.265 ;
        RECT 500.660 103.260 500.955 110.085 ;
        RECT 501.790 102.720 502.090 109.530 ;
        RECT 502.580 103.315 502.890 113.355 ;
        RECT 511.770 111.600 512.150 111.980 ;
        RECT 503.375 103.245 503.675 110.075 ;
        RECT 504.500 102.630 504.800 109.570 ;
        RECT 505.950 102.505 506.230 105.540 ;
        RECT 506.710 103.205 506.990 109.565 ;
        RECT 507.560 103.205 507.860 110.025 ;
        RECT 508.700 102.460 509.000 109.615 ;
        RECT 509.345 106.650 509.725 107.030 ;
        RECT 509.345 104.595 509.725 104.975 ;
        RECT 511.195 104.475 511.510 108.800 ;
        RECT 511.805 106.550 512.085 108.080 ;
        RECT 512.375 103.235 512.675 110.275 ;
        RECT 513.495 102.630 513.795 109.560 ;
        RECT 514.150 103.990 514.450 108.050 ;
        RECT 514.805 103.230 515.105 109.580 ;
        RECT 511.670 101.425 512.050 101.805 ;
        RECT 515.400 101.020 515.690 110.265 ;
        RECT 516.120 103.260 516.415 110.085 ;
        RECT 517.250 102.720 517.550 109.530 ;
        RECT 518.040 103.315 518.350 112.050 ;
        RECT 518.835 103.245 519.135 110.075 ;
        RECT 519.960 102.630 520.260 109.570 ;
        RECT 520.640 103.975 520.920 108.065 ;
        RECT 521.410 102.505 521.690 105.540 ;
        RECT 522.170 103.205 522.450 109.565 ;
        RECT 523.020 103.205 523.320 110.025 ;
        RECT 524.160 102.460 524.460 109.615 ;
        RECT 526.365 108.385 526.740 116.585 ;
        RECT 528.110 107.580 528.410 118.575 ;
        RECT 529.200 106.540 529.580 116.795 ;
        RECT 530.070 104.385 530.505 117.960 ;
        RECT 585.925 117.240 586.440 127.290 ;
        RECT 587.610 115.885 588.195 126.665 ;
        RECT 589.155 124.150 589.510 138.205 ;
        RECT 652.500 137.575 652.950 147.690 ;
        RECT 590.780 124.955 591.140 136.605 ;
        RECT 653.665 136.035 654.150 144.790 ;
        RECT 660.270 135.410 660.675 146.940 ;
        RECT 662.345 137.310 662.735 148.410 ;
        RECT 665.615 140.885 665.970 151.970 ;
        RECT 669.360 150.610 669.650 152.670 ;
        RECT 672.130 151.210 672.630 154.260 ;
        RECT 677.100 151.120 677.510 154.215 ;
        RECT 676.140 149.460 676.450 149.490 ;
        RECT 666.940 145.740 667.410 148.730 ;
        RECT 669.290 142.755 669.605 145.125 ;
        RECT 670.910 144.800 671.330 148.765 ;
        RECT 667.575 140.045 667.955 141.420 ;
        RECT 670.015 139.015 670.360 141.475 ;
        RECT 671.650 140.695 671.975 143.460 ;
        RECT 672.635 142.730 673.040 146.060 ;
        RECT 676.140 143.360 676.455 149.460 ;
        RECT 677.285 139.755 677.655 148.855 ;
        RECT 678.230 140.820 678.520 152.655 ;
        RECT 681.680 151.095 682.090 154.190 ;
        RECT 686.135 150.550 686.445 153.065 ;
        RECT 690.385 152.250 690.765 152.630 ;
        RECT 692.515 152.250 692.895 152.630 ;
        RECT 679.125 143.315 679.455 149.510 ;
        RECT 682.030 142.785 682.485 146.060 ;
        RECT 684.390 144.800 684.935 148.740 ;
        RECT 688.445 145.740 688.880 148.750 ;
        RECT 683.585 140.695 683.910 143.460 ;
        RECT 686.100 142.790 686.515 145.180 ;
        RECT 689.640 141.365 689.970 152.060 ;
        RECT 691.075 145.700 691.460 151.485 ;
        RECT 687.830 139.960 688.165 141.310 ;
        RECT 691.435 140.945 691.860 145.220 ;
        RECT 693.135 142.710 693.435 149.750 ;
        RECT 694.255 142.105 694.555 149.035 ;
        RECT 695.565 142.705 695.865 149.055 ;
        RECT 690.095 140.035 690.475 140.415 ;
        RECT 692.290 140.020 692.670 140.400 ;
        RECT 696.160 139.960 696.450 149.740 ;
        RECT 696.880 142.735 697.175 149.560 ;
        RECT 698.010 142.195 698.310 149.005 ;
        RECT 698.800 142.790 699.110 152.830 ;
        RECT 707.990 151.075 708.370 151.455 ;
        RECT 699.595 142.720 699.895 149.550 ;
        RECT 700.720 142.105 701.020 149.045 ;
        RECT 702.170 141.980 702.450 145.015 ;
        RECT 702.930 142.680 703.210 149.040 ;
        RECT 703.780 142.680 704.080 149.500 ;
        RECT 704.920 141.935 705.220 149.090 ;
        RECT 705.565 146.125 705.945 146.505 ;
        RECT 705.565 144.070 705.945 144.450 ;
        RECT 707.415 143.950 707.730 148.275 ;
        RECT 708.025 146.025 708.305 147.555 ;
        RECT 708.595 142.710 708.895 149.750 ;
        RECT 709.715 142.105 710.015 149.035 ;
        RECT 710.370 143.465 710.670 147.525 ;
        RECT 711.025 142.705 711.325 149.055 ;
        RECT 707.890 140.900 708.270 141.280 ;
        RECT 711.620 140.495 711.910 149.740 ;
        RECT 712.340 142.735 712.635 149.560 ;
        RECT 713.470 142.195 713.770 149.005 ;
        RECT 714.260 142.790 714.570 151.525 ;
        RECT 715.055 142.720 715.355 149.550 ;
        RECT 716.180 142.105 716.480 149.045 ;
        RECT 716.860 143.450 717.140 147.540 ;
        RECT 717.630 141.980 717.910 145.015 ;
        RECT 718.390 142.680 718.670 149.040 ;
        RECT 719.240 142.680 719.540 149.500 ;
        RECT 720.380 141.935 720.680 149.090 ;
        RECT 722.420 147.830 722.795 156.030 ;
        RECT 724.165 147.025 724.465 158.020 ;
        RECT 725.565 145.985 725.945 156.240 ;
        RECT 726.435 143.830 726.870 157.405 ;
        RECT 782.140 156.650 782.655 166.700 ;
        RECT 790.850 166.235 791.230 166.615 ;
        RECT 783.825 155.295 784.410 166.075 ;
        RECT 790.815 165.565 791.195 165.945 ;
        RECT 791.530 162.490 791.830 169.530 ;
        RECT 792.650 161.885 792.950 168.815 ;
        RECT 793.305 163.245 793.605 167.305 ;
        RECT 793.960 162.485 794.260 168.835 ;
        RECT 794.555 164.360 794.875 169.520 ;
        RECT 795.275 162.515 795.570 169.340 ;
        RECT 796.405 161.975 796.705 168.785 ;
        RECT 797.195 162.570 797.505 168.760 ;
        RECT 797.990 162.500 798.290 169.330 ;
        RECT 799.115 161.885 799.415 168.825 ;
        RECT 799.795 163.230 800.075 167.320 ;
        RECT 800.565 161.760 800.845 164.795 ;
        RECT 801.325 162.460 801.630 168.820 ;
        RECT 802.175 162.460 802.475 169.280 ;
        RECT 803.315 161.715 803.615 168.870 ;
        RECT 803.980 167.670 804.360 168.050 ;
        RECT 806.250 167.670 806.630 168.075 ;
        RECT 803.985 166.920 804.365 167.300 ;
        RECT 806.255 166.920 806.635 167.325 ;
        RECT 803.985 165.905 804.365 166.285 ;
        RECT 805.770 164.485 806.090 166.615 ;
        RECT 804.200 161.195 804.580 164.215 ;
        RECT 806.380 163.645 806.660 166.050 ;
        RECT 806.990 162.490 807.290 169.530 ;
        RECT 808.110 161.885 808.410 168.815 ;
        RECT 808.765 163.245 809.065 167.305 ;
        RECT 809.420 162.485 809.720 168.835 ;
        RECT 810.015 164.360 810.340 169.520 ;
        RECT 810.735 162.515 811.030 169.340 ;
        RECT 811.865 161.975 812.165 168.785 ;
        RECT 812.655 162.570 812.965 168.760 ;
        RECT 813.450 162.500 813.750 169.330 ;
        RECT 814.575 161.885 814.875 168.825 ;
        RECT 815.255 163.230 815.535 167.320 ;
        RECT 816.025 161.760 816.305 164.795 ;
        RECT 816.785 162.460 817.105 168.820 ;
        RECT 817.635 162.460 817.935 169.280 ;
        RECT 818.775 161.715 819.075 168.870 ;
        RECT 819.715 167.670 820.075 169.500 ;
        RECT 819.410 163.860 819.790 164.240 ;
        RECT 820.115 159.745 820.475 166.305 ;
        RECT 821.255 164.495 821.580 166.360 ;
        RECT 821.895 166.150 822.310 169.500 ;
        RECT 821.920 161.150 822.380 165.835 ;
        RECT 822.705 163.695 823.155 172.515 ;
        RECT 823.565 161.320 823.920 171.625 ;
        RECT 824.230 166.925 824.575 167.980 ;
        RECT 824.890 165.520 825.320 168.510 ;
        RECT 822.635 159.805 823.015 160.185 ;
        RECT 825.525 159.825 825.905 161.200 ;
        RECT 826.295 160.645 826.610 171.695 ;
        RECT 827.310 170.390 827.600 172.450 ;
        RECT 830.095 170.990 830.570 174.040 ;
        RECT 835.050 170.900 835.460 173.995 ;
        RECT 834.090 169.240 834.400 169.270 ;
        RECT 827.230 162.535 827.555 164.905 ;
        RECT 828.880 164.580 829.280 168.545 ;
        RECT 827.965 158.795 828.310 161.255 ;
        RECT 829.600 160.475 829.925 163.240 ;
        RECT 830.585 162.510 830.990 165.840 ;
        RECT 834.090 163.140 834.405 169.240 ;
        RECT 835.235 159.535 835.605 168.635 ;
        RECT 836.180 160.600 836.470 172.435 ;
        RECT 839.630 170.875 840.040 173.970 ;
        RECT 844.085 170.330 844.395 172.845 ;
        RECT 837.075 163.095 837.405 169.290 ;
        RECT 839.995 162.565 840.435 165.840 ;
        RECT 842.375 164.580 842.900 168.520 ;
        RECT 841.535 160.475 841.860 163.240 ;
        RECT 844.050 162.570 844.465 164.960 ;
        RECT 845.080 161.130 845.395 171.815 ;
        RECT 846.410 165.520 846.895 168.530 ;
        RECT 847.590 161.145 847.920 171.840 ;
        RECT 845.780 159.740 846.115 161.090 ;
        RECT 757.325 140.990 757.640 152.040 ;
        RECT 761.160 151.335 761.560 154.385 ;
        RECT 766.080 151.245 766.490 154.340 ;
        RECT 770.660 151.220 771.070 154.315 ;
        RECT 758.995 139.140 759.340 141.600 ;
        RECT 776.110 141.475 776.425 152.160 ;
        RECT 781.295 144.265 781.745 148.425 ;
        RECT 782.995 147.245 783.520 147.685 ;
        RECT 594.620 128.270 595.000 128.650 ;
        RECT 594.610 127.520 594.990 127.900 ;
        RECT 594.655 126.835 595.035 127.215 ;
        RECT 594.620 126.165 595.000 126.545 ;
        RECT 595.335 123.090 595.635 130.130 ;
        RECT 596.455 122.485 596.755 129.415 ;
        RECT 597.110 123.845 597.410 127.905 ;
        RECT 597.765 123.085 598.065 129.435 ;
        RECT 598.360 124.960 598.680 130.120 ;
        RECT 599.080 123.115 599.375 129.940 ;
        RECT 600.210 122.575 600.510 129.385 ;
        RECT 601.000 123.170 601.310 129.360 ;
        RECT 601.795 123.100 602.095 129.930 ;
        RECT 602.920 122.485 603.220 129.425 ;
        RECT 603.600 123.830 603.880 127.920 ;
        RECT 604.370 122.360 604.650 125.395 ;
        RECT 605.130 123.060 605.435 129.420 ;
        RECT 605.980 123.060 606.280 129.880 ;
        RECT 607.120 122.315 607.420 129.470 ;
        RECT 607.785 128.270 608.165 128.650 ;
        RECT 610.055 128.270 610.435 128.675 ;
        RECT 607.790 127.520 608.170 127.900 ;
        RECT 610.060 127.520 610.440 127.925 ;
        RECT 607.790 126.505 608.170 126.885 ;
        RECT 609.575 125.085 609.895 127.215 ;
        RECT 608.005 121.795 608.385 124.815 ;
        RECT 610.185 124.245 610.465 126.650 ;
        RECT 610.795 123.090 611.095 130.130 ;
        RECT 611.915 122.485 612.215 129.415 ;
        RECT 612.570 123.845 612.870 127.905 ;
        RECT 613.225 123.085 613.525 129.435 ;
        RECT 613.820 124.960 614.145 130.120 ;
        RECT 614.540 123.115 614.835 129.940 ;
        RECT 615.670 122.575 615.970 129.385 ;
        RECT 616.460 123.170 616.770 129.360 ;
        RECT 617.255 123.100 617.555 129.930 ;
        RECT 618.380 122.485 618.680 129.425 ;
        RECT 619.060 123.830 619.340 127.920 ;
        RECT 619.830 122.360 620.110 125.395 ;
        RECT 620.590 123.060 620.910 129.420 ;
        RECT 621.440 123.060 621.740 129.880 ;
        RECT 622.580 122.315 622.880 129.470 ;
        RECT 623.520 128.270 623.880 130.100 ;
        RECT 623.215 124.460 623.595 124.840 ;
        RECT 623.920 120.345 624.280 126.905 ;
        RECT 625.060 125.095 625.385 126.960 ;
        RECT 625.700 126.750 626.115 130.100 ;
        RECT 625.725 121.750 626.185 126.435 ;
        RECT 626.510 124.295 626.960 133.115 ;
        RECT 627.370 121.920 627.725 132.225 ;
        RECT 628.035 127.525 628.380 128.580 ;
        RECT 628.695 126.120 629.125 129.110 ;
        RECT 626.440 120.405 626.820 120.785 ;
        RECT 629.330 120.425 629.710 121.800 ;
        RECT 630.100 121.245 630.415 132.295 ;
        RECT 631.115 130.990 631.405 133.050 ;
        RECT 633.900 131.590 634.375 134.640 ;
        RECT 638.855 131.500 639.265 134.595 ;
        RECT 637.895 129.840 638.205 129.870 ;
        RECT 631.035 123.135 631.360 125.505 ;
        RECT 632.685 125.180 633.085 129.145 ;
        RECT 631.770 119.395 632.115 121.855 ;
        RECT 633.405 121.075 633.730 123.840 ;
        RECT 634.390 123.110 634.795 126.440 ;
        RECT 637.895 123.740 638.210 129.840 ;
        RECT 639.040 120.135 639.410 129.235 ;
        RECT 639.985 121.200 640.275 133.035 ;
        RECT 643.435 131.475 643.845 134.570 ;
        RECT 647.890 130.930 648.200 133.445 ;
        RECT 640.880 123.695 641.210 129.890 ;
        RECT 643.800 123.165 644.240 126.440 ;
        RECT 646.180 125.180 646.705 129.120 ;
        RECT 645.340 121.075 645.665 123.840 ;
        RECT 647.855 123.170 648.270 125.560 ;
        RECT 648.885 121.730 649.200 132.415 ;
        RECT 650.215 126.120 650.700 129.130 ;
        RECT 651.395 121.745 651.725 132.440 ;
        RECT 649.585 120.340 649.920 121.690 ;
        RECT 560.950 101.410 561.265 112.460 ;
        RECT 564.785 111.755 565.185 114.805 ;
        RECT 569.705 111.665 570.115 114.760 ;
        RECT 574.285 111.640 574.695 114.735 ;
        RECT 562.620 99.560 562.965 102.020 ;
        RECT 579.735 101.895 580.050 112.580 ;
        RECT 584.920 104.685 585.370 108.845 ;
        RECT 586.620 107.665 587.145 108.105 ;
        RECT 397.920 88.685 398.300 89.065 ;
        RECT 397.910 87.935 398.290 88.315 ;
        RECT 397.955 87.250 398.335 87.630 ;
        RECT 397.920 86.580 398.300 86.960 ;
        RECT 398.635 83.505 398.935 90.545 ;
        RECT 399.755 82.900 400.055 89.830 ;
        RECT 400.410 84.260 400.710 88.320 ;
        RECT 401.065 83.500 401.365 89.850 ;
        RECT 401.660 85.375 401.980 90.535 ;
        RECT 402.380 83.530 402.675 90.355 ;
        RECT 403.510 82.990 403.810 89.800 ;
        RECT 404.300 83.585 404.610 89.775 ;
        RECT 405.095 83.515 405.395 90.345 ;
        RECT 406.220 82.900 406.520 89.840 ;
        RECT 406.900 84.245 407.180 88.335 ;
        RECT 407.670 82.775 407.950 85.810 ;
        RECT 408.430 83.475 408.735 89.835 ;
        RECT 409.280 83.475 409.580 90.295 ;
        RECT 410.420 82.730 410.720 89.885 ;
        RECT 411.085 88.685 411.465 89.065 ;
        RECT 413.355 88.685 413.735 89.090 ;
        RECT 411.090 87.935 411.470 88.315 ;
        RECT 413.360 87.935 413.740 88.340 ;
        RECT 411.090 86.920 411.470 87.300 ;
        RECT 412.875 85.500 413.195 87.630 ;
        RECT 411.305 82.210 411.685 85.230 ;
        RECT 413.485 84.660 413.765 87.065 ;
        RECT 414.095 83.505 414.395 90.545 ;
        RECT 415.215 82.900 415.515 89.830 ;
        RECT 415.870 84.260 416.170 88.320 ;
        RECT 416.525 83.500 416.825 89.850 ;
        RECT 417.120 85.375 417.445 90.535 ;
        RECT 417.840 83.530 418.135 90.355 ;
        RECT 418.970 82.990 419.270 89.800 ;
        RECT 419.760 83.585 420.070 89.775 ;
        RECT 420.555 83.515 420.855 90.345 ;
        RECT 421.680 82.900 421.980 89.840 ;
        RECT 422.360 84.245 422.640 88.335 ;
        RECT 423.130 82.775 423.410 85.810 ;
        RECT 423.890 83.475 424.210 89.835 ;
        RECT 424.740 83.475 425.040 90.295 ;
        RECT 425.880 82.730 426.180 89.885 ;
        RECT 426.820 88.685 427.180 90.515 ;
        RECT 426.515 84.875 426.895 85.255 ;
        RECT 427.220 80.760 427.580 87.320 ;
        RECT 428.360 85.510 428.685 87.375 ;
        RECT 429.000 87.165 429.415 90.515 ;
        RECT 429.025 82.165 429.485 86.850 ;
        RECT 429.810 84.710 430.260 93.530 ;
        RECT 430.670 82.335 431.025 92.640 ;
        RECT 431.335 87.940 431.680 88.995 ;
        RECT 431.995 86.535 432.425 89.525 ;
        RECT 429.740 80.820 430.120 81.200 ;
        RECT 432.630 80.840 433.010 82.215 ;
        RECT 433.400 81.660 433.715 92.710 ;
        RECT 434.415 91.405 434.705 93.465 ;
        RECT 437.200 92.005 437.675 95.055 ;
        RECT 442.155 91.915 442.565 95.010 ;
        RECT 441.195 90.255 441.505 90.285 ;
        RECT 434.335 83.550 434.660 85.920 ;
        RECT 435.985 85.595 436.385 89.560 ;
        RECT 435.070 79.810 435.415 82.270 ;
        RECT 436.705 81.490 437.030 84.255 ;
        RECT 437.690 83.525 438.095 86.855 ;
        RECT 441.195 84.155 441.510 90.255 ;
        RECT 442.340 80.550 442.710 89.650 ;
        RECT 443.285 81.615 443.575 93.450 ;
        RECT 446.735 91.890 447.145 94.985 ;
        RECT 451.190 91.345 451.500 93.860 ;
        RECT 444.180 84.110 444.510 90.305 ;
        RECT 447.100 83.580 447.540 86.855 ;
        RECT 449.480 85.595 450.005 89.535 ;
        RECT 448.640 81.490 448.965 84.255 ;
        RECT 451.155 83.585 451.570 85.975 ;
        RECT 452.185 82.145 452.500 92.830 ;
        RECT 453.515 86.535 454.000 89.545 ;
        RECT 454.695 82.160 455.025 92.855 ;
        RECT 452.885 80.755 453.220 82.105 ;
        RECT 364.590 61.810 364.905 72.860 ;
        RECT 368.425 72.155 368.825 75.205 ;
        RECT 373.345 72.065 373.755 75.160 ;
        RECT 377.925 72.040 378.335 75.135 ;
        RECT 366.260 59.960 366.605 62.420 ;
        RECT 383.375 62.295 383.690 72.980 ;
        RECT 388.560 65.085 389.010 69.245 ;
        RECT 390.260 68.065 390.785 68.505 ;
        RECT 201.600 49.165 201.980 49.545 ;
        RECT 201.590 48.415 201.970 48.795 ;
        RECT 201.635 47.730 202.015 48.110 ;
        RECT 201.600 47.060 201.980 47.440 ;
        RECT 202.315 43.985 202.615 51.025 ;
        RECT 203.435 43.380 203.735 50.310 ;
        RECT 204.090 44.740 204.390 48.800 ;
        RECT 204.745 43.980 205.045 50.330 ;
        RECT 205.340 45.855 205.660 51.015 ;
        RECT 206.060 44.010 206.355 50.835 ;
        RECT 207.190 43.470 207.490 50.280 ;
        RECT 207.980 44.065 208.290 50.255 ;
        RECT 208.775 43.995 209.075 50.825 ;
        RECT 209.900 43.380 210.200 50.320 ;
        RECT 210.580 44.725 210.860 48.815 ;
        RECT 211.350 43.255 211.630 46.290 ;
        RECT 212.110 43.955 212.415 50.315 ;
        RECT 212.960 43.955 213.260 50.775 ;
        RECT 214.100 43.210 214.400 50.365 ;
        RECT 214.765 49.165 215.145 49.545 ;
        RECT 217.035 49.165 217.415 49.570 ;
        RECT 214.770 48.415 215.150 48.795 ;
        RECT 217.040 48.415 217.420 48.820 ;
        RECT 214.770 47.400 215.150 47.780 ;
        RECT 216.555 45.980 216.875 48.110 ;
        RECT 214.985 42.690 215.365 45.710 ;
        RECT 217.165 45.140 217.445 47.545 ;
        RECT 217.775 43.985 218.075 51.025 ;
        RECT 218.895 43.380 219.195 50.310 ;
        RECT 219.550 44.740 219.850 48.800 ;
        RECT 220.205 43.980 220.505 50.330 ;
        RECT 220.800 45.855 221.125 51.015 ;
        RECT 221.520 44.010 221.815 50.835 ;
        RECT 222.650 43.470 222.950 50.280 ;
        RECT 223.440 44.065 223.750 50.255 ;
        RECT 224.235 43.995 224.535 50.825 ;
        RECT 225.360 43.380 225.660 50.320 ;
        RECT 226.040 44.725 226.320 48.815 ;
        RECT 226.810 43.255 227.090 46.290 ;
        RECT 227.570 43.955 227.890 50.315 ;
        RECT 228.420 43.955 228.720 50.775 ;
        RECT 229.560 43.210 229.860 50.365 ;
        RECT 230.500 49.165 230.860 50.995 ;
        RECT 230.195 45.355 230.575 45.735 ;
        RECT 230.900 41.240 231.260 47.800 ;
        RECT 232.040 45.990 232.365 47.855 ;
        RECT 232.680 47.645 233.095 50.995 ;
        RECT 232.705 42.645 233.165 47.330 ;
        RECT 233.490 45.190 233.940 54.010 ;
        RECT 234.350 42.815 234.705 53.120 ;
        RECT 235.015 48.420 235.360 49.475 ;
        RECT 235.675 47.015 236.105 50.005 ;
        RECT 233.420 41.300 233.800 41.680 ;
        RECT 236.310 41.320 236.690 42.695 ;
        RECT 237.080 42.140 237.395 53.190 ;
        RECT 238.095 51.885 238.385 53.945 ;
        RECT 240.880 52.485 241.355 55.535 ;
        RECT 245.835 52.395 246.245 55.490 ;
        RECT 244.875 50.735 245.185 50.765 ;
        RECT 238.015 44.030 238.340 46.400 ;
        RECT 239.665 46.075 240.065 50.040 ;
        RECT 238.750 40.290 239.095 42.750 ;
        RECT 240.385 41.970 240.710 44.735 ;
        RECT 241.370 44.005 241.775 47.335 ;
        RECT 244.875 44.635 245.190 50.735 ;
        RECT 246.020 41.030 246.390 50.130 ;
        RECT 246.965 42.095 247.255 53.930 ;
        RECT 250.415 52.370 250.825 55.465 ;
        RECT 254.870 51.825 255.180 54.340 ;
        RECT 247.860 44.590 248.190 50.785 ;
        RECT 250.780 44.060 251.220 47.335 ;
        RECT 253.160 46.075 253.685 50.015 ;
        RECT 252.320 41.970 252.645 44.735 ;
        RECT 254.835 44.065 255.250 46.455 ;
        RECT 255.865 42.625 256.180 53.310 ;
        RECT 257.195 47.015 257.680 50.025 ;
        RECT 258.375 42.640 258.705 53.335 ;
        RECT 256.565 41.235 256.900 42.585 ;
        RECT 168.245 22.400 168.560 33.450 ;
        RECT 172.080 32.745 172.480 35.795 ;
        RECT 177.000 32.655 177.410 35.750 ;
        RECT 181.580 32.630 181.990 35.725 ;
        RECT 169.915 20.550 170.260 23.010 ;
        RECT 187.030 22.885 187.345 33.570 ;
        RECT 192.265 25.600 192.715 29.760 ;
        RECT 193.965 28.580 194.490 29.020 ;
        RECT 76.675 3.840 76.975 10.770 ;
        RECT 77.330 5.200 77.630 9.260 ;
        RECT 77.985 4.440 78.285 10.790 ;
        RECT 79.300 4.470 79.595 11.295 ;
        RECT 83.140 3.840 83.440 10.780 ;
        RECT 83.820 5.185 84.100 9.275 ;
        RECT 85.350 4.415 85.655 10.775 ;
        RECT 86.200 4.415 86.500 11.235 ;
        RECT 87.940 8.235 88.320 8.255 ;
        RECT 87.930 7.875 88.320 8.235 ;
        RECT 87.930 7.855 88.310 7.875 ;
        RECT 87.940 5.810 88.320 6.190 ;
        RECT 193.065 5.440 193.580 27.700 ;
        RECT 194.750 7.655 195.335 28.350 ;
        RECT 196.335 25.235 196.690 39.175 ;
        RECT 259.680 38.545 260.130 48.810 ;
        RECT 197.960 26.025 198.320 37.575 ;
        RECT 260.845 37.005 261.330 45.890 ;
        RECT 267.785 36.280 268.190 48.325 ;
        RECT 269.860 38.180 270.250 49.605 ;
        RECT 273.020 42.020 273.375 53.105 ;
        RECT 276.765 51.745 277.055 53.805 ;
        RECT 279.535 52.345 280.035 55.395 ;
        RECT 284.505 52.255 284.915 55.350 ;
        RECT 283.545 50.595 283.855 50.625 ;
        RECT 274.345 46.875 274.815 49.865 ;
        RECT 276.695 43.890 277.010 46.260 ;
        RECT 278.315 45.935 278.735 49.900 ;
        RECT 274.980 41.180 275.360 42.555 ;
        RECT 277.420 40.150 277.765 42.610 ;
        RECT 279.055 41.830 279.380 44.595 ;
        RECT 280.040 43.865 280.445 47.195 ;
        RECT 283.545 44.495 283.860 50.595 ;
        RECT 284.690 40.890 285.060 49.990 ;
        RECT 285.635 41.955 285.925 53.790 ;
        RECT 289.085 52.230 289.495 55.325 ;
        RECT 293.540 51.685 293.850 54.200 ;
        RECT 297.790 53.385 298.170 53.765 ;
        RECT 299.920 53.385 300.300 53.765 ;
        RECT 286.530 44.450 286.860 50.645 ;
        RECT 289.435 43.920 289.890 47.195 ;
        RECT 291.795 45.935 292.340 49.875 ;
        RECT 295.850 46.875 296.285 49.885 ;
        RECT 290.990 41.830 291.315 44.595 ;
        RECT 293.505 43.925 293.920 46.315 ;
        RECT 297.045 42.500 297.375 53.195 ;
        RECT 298.480 46.835 298.865 52.620 ;
        RECT 295.235 41.095 295.570 42.445 ;
        RECT 298.840 42.080 299.265 46.355 ;
        RECT 300.540 43.845 300.840 50.885 ;
        RECT 301.660 43.240 301.960 50.170 ;
        RECT 302.970 43.840 303.270 50.190 ;
        RECT 297.500 41.170 297.880 41.550 ;
        RECT 299.695 41.155 300.075 41.535 ;
        RECT 303.565 41.095 303.855 50.875 ;
        RECT 304.285 43.870 304.580 50.695 ;
        RECT 305.415 43.330 305.715 50.140 ;
        RECT 306.205 43.925 306.515 53.965 ;
        RECT 315.395 52.210 315.775 52.590 ;
        RECT 307.000 43.855 307.300 50.685 ;
        RECT 308.125 43.240 308.425 50.180 ;
        RECT 309.575 43.115 309.855 46.150 ;
        RECT 310.335 43.815 310.615 50.175 ;
        RECT 311.185 43.815 311.485 50.635 ;
        RECT 312.325 43.070 312.625 50.225 ;
        RECT 312.970 47.260 313.350 47.640 ;
        RECT 312.970 45.205 313.350 45.585 ;
        RECT 314.820 45.085 315.135 49.410 ;
        RECT 315.430 47.160 315.710 48.690 ;
        RECT 316.000 43.845 316.300 50.885 ;
        RECT 317.120 43.240 317.420 50.170 ;
        RECT 317.775 44.600 318.075 48.660 ;
        RECT 318.430 43.840 318.730 50.190 ;
        RECT 315.295 42.035 315.675 42.415 ;
        RECT 319.025 41.630 319.315 50.875 ;
        RECT 319.745 43.870 320.040 50.695 ;
        RECT 320.875 43.330 321.175 50.140 ;
        RECT 321.665 43.925 321.975 52.660 ;
        RECT 322.460 43.855 322.760 50.685 ;
        RECT 323.585 43.240 323.885 50.180 ;
        RECT 324.265 44.585 324.545 48.675 ;
        RECT 325.035 43.115 325.315 46.150 ;
        RECT 325.795 43.815 326.075 50.175 ;
        RECT 326.645 43.815 326.945 50.635 ;
        RECT 327.785 43.070 328.085 50.225 ;
        RECT 330.125 48.840 330.500 57.040 ;
        RECT 331.870 48.035 332.170 59.030 ;
        RECT 332.880 47.055 333.260 57.310 ;
        RECT 333.750 44.900 334.185 58.475 ;
        RECT 389.460 57.635 389.975 67.935 ;
        RECT 391.145 56.530 391.730 67.310 ;
        RECT 392.640 64.790 392.995 78.710 ;
        RECT 455.985 78.080 456.435 88.345 ;
        RECT 394.265 65.695 394.625 77.110 ;
        RECT 457.150 76.540 457.635 85.425 ;
        RECT 463.815 76.275 464.220 87.805 ;
        RECT 465.890 78.175 466.280 89.275 ;
        RECT 469.315 81.655 469.670 92.740 ;
        RECT 473.060 91.380 473.350 93.440 ;
        RECT 475.830 91.980 476.330 95.030 ;
        RECT 480.800 91.890 481.210 94.985 ;
        RECT 479.840 90.230 480.150 90.260 ;
        RECT 470.640 86.510 471.110 89.500 ;
        RECT 472.990 83.525 473.305 85.895 ;
        RECT 474.610 85.570 475.030 89.535 ;
        RECT 471.275 80.815 471.655 82.190 ;
        RECT 473.715 79.785 474.060 82.245 ;
        RECT 475.350 81.465 475.675 84.230 ;
        RECT 476.335 83.500 476.740 86.830 ;
        RECT 479.840 84.130 480.155 90.230 ;
        RECT 480.985 80.525 481.355 89.625 ;
        RECT 481.930 81.590 482.220 93.425 ;
        RECT 485.380 91.865 485.790 94.960 ;
        RECT 489.835 91.320 490.145 93.835 ;
        RECT 494.085 93.020 494.465 93.400 ;
        RECT 496.215 93.020 496.595 93.400 ;
        RECT 482.825 84.085 483.155 90.280 ;
        RECT 485.730 83.555 486.185 86.830 ;
        RECT 488.090 85.570 488.635 89.510 ;
        RECT 492.145 86.510 492.580 89.520 ;
        RECT 487.285 81.465 487.610 84.230 ;
        RECT 489.800 83.560 490.215 85.950 ;
        RECT 493.340 82.135 493.670 92.830 ;
        RECT 494.775 86.470 495.160 92.255 ;
        RECT 491.530 80.730 491.865 82.080 ;
        RECT 495.135 81.715 495.560 85.990 ;
        RECT 496.835 83.480 497.135 90.520 ;
        RECT 497.955 82.875 498.255 89.805 ;
        RECT 499.265 83.475 499.565 89.825 ;
        RECT 493.795 80.805 494.175 81.185 ;
        RECT 495.990 80.790 496.370 81.170 ;
        RECT 499.860 80.730 500.150 90.510 ;
        RECT 500.580 83.505 500.875 90.330 ;
        RECT 501.710 82.965 502.010 89.775 ;
        RECT 502.500 83.560 502.810 93.600 ;
        RECT 511.690 91.845 512.070 92.225 ;
        RECT 503.295 83.490 503.595 90.320 ;
        RECT 504.420 82.875 504.720 89.815 ;
        RECT 505.870 82.750 506.150 85.785 ;
        RECT 506.630 83.450 506.910 89.810 ;
        RECT 507.480 83.450 507.780 90.270 ;
        RECT 508.620 82.705 508.920 89.860 ;
        RECT 509.265 86.895 509.645 87.275 ;
        RECT 509.265 84.840 509.645 85.220 ;
        RECT 511.115 84.720 511.430 89.045 ;
        RECT 511.725 86.795 512.005 88.325 ;
        RECT 512.295 83.480 512.595 90.520 ;
        RECT 513.415 82.875 513.715 89.805 ;
        RECT 514.070 84.235 514.370 88.295 ;
        RECT 514.725 83.475 515.025 89.825 ;
        RECT 511.590 81.670 511.970 82.050 ;
        RECT 515.320 81.265 515.610 90.510 ;
        RECT 516.040 83.505 516.335 90.330 ;
        RECT 517.170 82.965 517.470 89.775 ;
        RECT 517.960 83.560 518.270 92.295 ;
        RECT 518.755 83.490 519.055 90.320 ;
        RECT 519.880 82.875 520.180 89.815 ;
        RECT 520.560 84.220 520.840 88.310 ;
        RECT 521.330 82.750 521.610 85.785 ;
        RECT 522.090 83.450 522.370 89.810 ;
        RECT 522.940 83.450 523.240 90.270 ;
        RECT 524.080 82.705 524.380 89.860 ;
        RECT 526.365 88.565 526.740 96.850 ;
        RECT 528.110 87.845 528.410 98.840 ;
        RECT 529.200 86.785 529.580 97.040 ;
        RECT 530.070 84.630 530.505 98.205 ;
        RECT 585.775 97.405 586.290 107.455 ;
        RECT 587.460 96.050 588.045 106.830 ;
        RECT 589.365 104.375 589.720 118.165 ;
        RECT 652.710 117.535 653.160 128.035 ;
        RECT 590.990 105.230 591.350 116.565 ;
        RECT 653.875 115.995 654.360 125.235 ;
        RECT 660.290 115.750 660.695 127.280 ;
        RECT 662.365 117.650 662.755 128.750 ;
        RECT 665.770 121.240 666.125 132.325 ;
        RECT 669.515 130.965 669.805 133.025 ;
        RECT 672.285 131.565 672.785 134.615 ;
        RECT 677.255 131.475 677.665 134.570 ;
        RECT 676.295 129.815 676.605 129.845 ;
        RECT 667.095 126.095 667.565 129.085 ;
        RECT 669.445 123.110 669.760 125.480 ;
        RECT 671.065 125.155 671.485 129.120 ;
        RECT 667.730 120.400 668.110 121.775 ;
        RECT 670.170 119.370 670.515 121.830 ;
        RECT 671.805 121.050 672.130 123.815 ;
        RECT 672.790 123.085 673.195 126.415 ;
        RECT 676.295 123.715 676.610 129.815 ;
        RECT 677.440 120.110 677.810 129.210 ;
        RECT 678.385 121.175 678.675 133.010 ;
        RECT 681.835 131.450 682.245 134.545 ;
        RECT 686.290 130.905 686.600 133.420 ;
        RECT 690.540 132.605 690.920 132.985 ;
        RECT 692.670 132.605 693.050 132.985 ;
        RECT 679.280 123.670 679.610 129.865 ;
        RECT 682.185 123.140 682.640 126.415 ;
        RECT 684.545 125.155 685.090 129.095 ;
        RECT 688.600 126.095 689.035 129.105 ;
        RECT 683.740 121.050 684.065 123.815 ;
        RECT 686.255 123.145 686.670 125.535 ;
        RECT 689.795 121.720 690.125 132.415 ;
        RECT 691.230 126.055 691.615 131.840 ;
        RECT 687.985 120.315 688.320 121.665 ;
        RECT 691.590 121.300 692.015 125.575 ;
        RECT 693.290 123.065 693.590 130.105 ;
        RECT 694.410 122.460 694.710 129.390 ;
        RECT 695.720 123.060 696.020 129.410 ;
        RECT 690.250 120.390 690.630 120.770 ;
        RECT 692.445 120.375 692.825 120.755 ;
        RECT 696.315 120.315 696.605 130.095 ;
        RECT 697.035 123.090 697.330 129.915 ;
        RECT 698.165 122.550 698.465 129.360 ;
        RECT 698.955 123.145 699.265 133.185 ;
        RECT 708.145 131.430 708.525 131.810 ;
        RECT 699.750 123.075 700.050 129.905 ;
        RECT 700.875 122.460 701.175 129.400 ;
        RECT 702.325 122.335 702.605 125.370 ;
        RECT 703.085 123.035 703.365 129.395 ;
        RECT 703.935 123.035 704.235 129.855 ;
        RECT 705.075 122.290 705.375 129.445 ;
        RECT 705.720 126.480 706.100 126.860 ;
        RECT 705.720 124.425 706.100 124.805 ;
        RECT 707.570 124.305 707.885 128.630 ;
        RECT 708.180 126.380 708.460 127.910 ;
        RECT 708.750 123.065 709.050 130.105 ;
        RECT 709.870 122.460 710.170 129.390 ;
        RECT 710.525 123.820 710.825 127.880 ;
        RECT 711.180 123.060 711.480 129.410 ;
        RECT 708.045 121.255 708.425 121.635 ;
        RECT 711.775 120.850 712.065 130.095 ;
        RECT 712.495 123.090 712.790 129.915 ;
        RECT 713.625 122.550 713.925 129.360 ;
        RECT 714.415 123.145 714.725 131.880 ;
        RECT 715.210 123.075 715.510 129.905 ;
        RECT 716.335 122.460 716.635 129.400 ;
        RECT 717.015 123.805 717.295 127.895 ;
        RECT 717.785 122.335 718.065 125.370 ;
        RECT 718.545 123.035 718.825 129.395 ;
        RECT 719.395 123.035 719.695 129.855 ;
        RECT 720.535 122.290 720.835 129.445 ;
        RECT 722.720 128.080 723.095 136.280 ;
        RECT 724.465 127.275 724.765 138.270 ;
        RECT 725.565 126.340 725.945 136.595 ;
        RECT 726.435 124.185 726.870 137.760 ;
        RECT 782.140 136.960 782.655 147.010 ;
        RECT 783.825 135.605 784.410 146.385 ;
        RECT 785.495 143.915 785.850 157.705 ;
        RECT 848.840 157.075 849.290 167.340 ;
        RECT 787.120 144.770 787.480 156.105 ;
        RECT 850.005 155.535 850.490 164.420 ;
        RECT 856.310 155.160 856.715 166.690 ;
        RECT 858.385 157.060 858.775 168.160 ;
        RECT 862.155 160.610 862.510 171.695 ;
        RECT 865.900 170.335 866.190 172.395 ;
        RECT 868.670 170.935 869.170 173.985 ;
        RECT 873.640 170.845 874.050 173.940 ;
        RECT 872.680 169.185 872.990 169.215 ;
        RECT 863.480 165.465 863.950 168.455 ;
        RECT 865.830 162.480 866.145 164.850 ;
        RECT 867.450 164.525 867.870 168.490 ;
        RECT 864.115 159.770 864.495 161.145 ;
        RECT 866.555 158.740 866.900 161.200 ;
        RECT 868.190 160.420 868.515 163.185 ;
        RECT 869.175 162.455 869.580 165.785 ;
        RECT 872.680 163.085 872.995 169.185 ;
        RECT 873.825 159.480 874.195 168.580 ;
        RECT 874.770 160.545 875.060 172.380 ;
        RECT 878.220 170.820 878.630 173.915 ;
        RECT 882.675 170.275 882.985 172.790 ;
        RECT 886.925 171.975 887.305 172.355 ;
        RECT 889.055 171.975 889.435 172.355 ;
        RECT 875.665 163.040 875.995 169.235 ;
        RECT 878.570 162.510 879.025 165.785 ;
        RECT 880.930 164.525 881.475 168.465 ;
        RECT 884.985 165.465 885.420 168.475 ;
        RECT 880.125 160.420 880.450 163.185 ;
        RECT 882.640 162.515 883.055 164.905 ;
        RECT 886.180 161.090 886.510 171.785 ;
        RECT 887.615 165.425 888.000 171.210 ;
        RECT 884.370 159.685 884.705 161.035 ;
        RECT 887.975 160.670 888.400 164.945 ;
        RECT 889.675 162.435 889.975 169.475 ;
        RECT 890.795 161.830 891.095 168.760 ;
        RECT 892.105 162.430 892.405 168.780 ;
        RECT 886.635 159.760 887.015 160.140 ;
        RECT 888.830 159.745 889.210 160.125 ;
        RECT 892.700 159.685 892.990 169.465 ;
        RECT 893.420 162.460 893.715 169.285 ;
        RECT 894.550 161.920 894.850 168.730 ;
        RECT 895.340 162.515 895.650 172.555 ;
        RECT 904.530 170.800 904.910 171.180 ;
        RECT 896.135 162.445 896.435 169.275 ;
        RECT 897.260 161.830 897.560 168.770 ;
        RECT 898.710 161.705 898.990 164.740 ;
        RECT 899.470 162.405 899.750 168.765 ;
        RECT 900.320 162.405 900.620 169.225 ;
        RECT 901.460 161.660 901.760 168.815 ;
        RECT 902.105 165.850 902.485 166.230 ;
        RECT 902.105 163.795 902.485 164.175 ;
        RECT 903.955 163.675 904.270 168.000 ;
        RECT 904.565 165.750 904.845 167.280 ;
        RECT 905.135 162.435 905.435 169.475 ;
        RECT 906.910 163.190 907.210 167.250 ;
        RECT 904.430 160.625 904.810 161.005 ;
        RECT 908.160 160.220 908.450 169.465 ;
        RECT 910.010 161.920 910.310 168.730 ;
        RECT 910.800 162.515 911.110 171.250 ;
        RECT 911.595 162.445 911.895 169.275 ;
        RECT 913.400 163.175 913.680 167.265 ;
        RECT 914.170 161.705 914.450 164.740 ;
        RECT 916.920 161.660 917.220 168.815 ;
        RECT 953.795 160.690 954.110 171.740 ;
        RECT 957.630 171.035 958.030 174.085 ;
        RECT 962.550 170.945 962.960 174.040 ;
        RECT 967.130 170.920 967.540 174.015 ;
        RECT 955.465 158.840 955.810 161.300 ;
        RECT 972.580 161.175 972.895 171.860 ;
        RECT 977.765 163.965 978.215 168.125 ;
        RECT 987.155 167.670 987.535 168.050 ;
        RECT 979.465 166.945 979.990 167.385 ;
        RECT 987.145 166.920 987.525 167.300 ;
        RECT 790.770 147.980 791.150 148.360 ;
        RECT 790.760 147.230 791.140 147.610 ;
        RECT 790.805 146.545 791.185 146.925 ;
        RECT 790.770 145.875 791.150 146.255 ;
        RECT 791.485 142.800 791.785 149.840 ;
        RECT 792.605 142.195 792.905 149.125 ;
        RECT 793.260 143.555 793.560 147.615 ;
        RECT 793.915 142.795 794.215 149.145 ;
        RECT 794.510 144.670 794.830 149.830 ;
        RECT 795.230 142.825 795.525 149.650 ;
        RECT 796.360 142.285 796.660 149.095 ;
        RECT 797.150 142.880 797.460 149.070 ;
        RECT 797.945 142.810 798.245 149.640 ;
        RECT 799.070 142.195 799.370 149.135 ;
        RECT 799.750 143.540 800.030 147.630 ;
        RECT 800.520 142.070 800.800 145.105 ;
        RECT 801.280 142.770 801.585 149.130 ;
        RECT 802.130 142.770 802.430 149.590 ;
        RECT 803.270 142.025 803.570 149.180 ;
        RECT 803.935 147.980 804.315 148.360 ;
        RECT 806.205 147.980 806.585 148.385 ;
        RECT 803.940 147.230 804.320 147.610 ;
        RECT 806.210 147.230 806.590 147.635 ;
        RECT 803.940 146.215 804.320 146.595 ;
        RECT 805.725 144.795 806.045 146.925 ;
        RECT 804.155 141.505 804.535 144.525 ;
        RECT 806.335 143.955 806.615 146.360 ;
        RECT 806.945 142.800 807.245 149.840 ;
        RECT 808.065 142.195 808.365 149.125 ;
        RECT 808.720 143.555 809.020 147.615 ;
        RECT 809.375 142.795 809.675 149.145 ;
        RECT 809.970 144.670 810.295 149.830 ;
        RECT 810.690 142.825 810.985 149.650 ;
        RECT 811.820 142.285 812.120 149.095 ;
        RECT 812.610 142.880 812.920 149.070 ;
        RECT 813.405 142.810 813.705 149.640 ;
        RECT 814.530 142.195 814.830 149.135 ;
        RECT 815.210 143.540 815.490 147.630 ;
        RECT 815.980 142.070 816.260 145.105 ;
        RECT 816.740 142.770 817.060 149.130 ;
        RECT 817.590 142.770 817.890 149.590 ;
        RECT 818.730 142.025 819.030 149.180 ;
        RECT 819.670 147.980 820.030 149.810 ;
        RECT 819.365 144.170 819.745 144.550 ;
        RECT 820.070 140.055 820.430 146.615 ;
        RECT 821.210 144.805 821.535 146.670 ;
        RECT 821.850 146.460 822.265 149.810 ;
        RECT 821.875 141.460 822.335 146.145 ;
        RECT 822.660 144.005 823.110 152.825 ;
        RECT 823.520 141.630 823.875 151.935 ;
        RECT 824.185 147.235 824.530 148.290 ;
        RECT 824.845 145.830 825.275 148.820 ;
        RECT 822.590 140.115 822.970 140.495 ;
        RECT 825.480 140.135 825.860 141.510 ;
        RECT 826.250 140.955 826.565 152.005 ;
        RECT 827.265 150.700 827.555 152.760 ;
        RECT 830.050 151.300 830.525 154.350 ;
        RECT 835.005 151.210 835.415 154.305 ;
        RECT 834.045 149.550 834.355 149.580 ;
        RECT 827.185 142.845 827.510 145.215 ;
        RECT 828.835 144.890 829.235 148.855 ;
        RECT 827.920 139.105 828.265 141.565 ;
        RECT 829.555 140.785 829.880 143.550 ;
        RECT 830.540 142.820 830.945 146.150 ;
        RECT 834.045 143.450 834.360 149.550 ;
        RECT 835.190 139.845 835.560 148.945 ;
        RECT 836.135 140.910 836.425 152.745 ;
        RECT 839.585 151.185 839.995 154.280 ;
        RECT 844.040 150.640 844.350 153.155 ;
        RECT 837.030 143.405 837.360 149.600 ;
        RECT 839.950 142.875 840.390 146.150 ;
        RECT 842.330 144.890 842.855 148.830 ;
        RECT 841.490 140.785 841.815 143.550 ;
        RECT 844.005 142.880 844.420 145.270 ;
        RECT 845.035 141.440 845.350 152.125 ;
        RECT 846.365 145.830 846.850 148.840 ;
        RECT 847.545 141.455 847.875 152.150 ;
        RECT 845.735 140.050 846.070 141.400 ;
        RECT 757.385 121.185 757.700 132.235 ;
        RECT 761.220 131.530 761.620 134.580 ;
        RECT 766.140 131.440 766.550 134.535 ;
        RECT 770.720 131.415 771.130 134.510 ;
        RECT 759.055 119.335 759.400 121.795 ;
        RECT 776.170 121.670 776.485 132.355 ;
        RECT 781.355 124.460 781.805 128.620 ;
        RECT 783.055 127.440 783.580 127.880 ;
        RECT 594.425 108.430 594.805 108.810 ;
        RECT 594.415 107.680 594.795 108.060 ;
        RECT 594.460 106.995 594.840 107.375 ;
        RECT 594.425 106.325 594.805 106.705 ;
        RECT 595.140 103.250 595.440 110.290 ;
        RECT 596.260 102.645 596.560 109.575 ;
        RECT 596.915 104.005 597.215 108.065 ;
        RECT 597.570 103.245 597.870 109.595 ;
        RECT 598.165 105.120 598.485 110.280 ;
        RECT 598.885 103.275 599.180 110.100 ;
        RECT 600.015 102.735 600.315 109.545 ;
        RECT 600.805 103.330 601.115 109.520 ;
        RECT 601.600 103.260 601.900 110.090 ;
        RECT 602.725 102.645 603.025 109.585 ;
        RECT 603.405 103.990 603.685 108.080 ;
        RECT 604.175 102.520 604.455 105.555 ;
        RECT 604.935 103.220 605.240 109.580 ;
        RECT 605.785 103.220 606.085 110.040 ;
        RECT 606.925 102.475 607.225 109.630 ;
        RECT 607.590 108.430 607.970 108.810 ;
        RECT 609.860 108.430 610.240 108.835 ;
        RECT 607.595 107.680 607.975 108.060 ;
        RECT 609.865 107.680 610.245 108.085 ;
        RECT 607.595 106.665 607.975 107.045 ;
        RECT 609.380 105.245 609.700 107.375 ;
        RECT 607.810 101.955 608.190 104.975 ;
        RECT 609.990 104.405 610.270 106.810 ;
        RECT 610.600 103.250 610.900 110.290 ;
        RECT 611.720 102.645 612.020 109.575 ;
        RECT 612.375 104.005 612.675 108.065 ;
        RECT 613.030 103.245 613.330 109.595 ;
        RECT 613.625 105.120 613.950 110.280 ;
        RECT 614.345 103.275 614.640 110.100 ;
        RECT 615.475 102.735 615.775 109.545 ;
        RECT 616.265 103.330 616.575 109.520 ;
        RECT 617.060 103.260 617.360 110.090 ;
        RECT 618.185 102.645 618.485 109.585 ;
        RECT 618.865 103.990 619.145 108.080 ;
        RECT 619.635 102.520 619.915 105.555 ;
        RECT 620.395 103.220 620.715 109.580 ;
        RECT 621.245 103.220 621.545 110.040 ;
        RECT 622.385 102.475 622.685 109.630 ;
        RECT 623.325 108.430 623.685 110.260 ;
        RECT 623.020 104.620 623.400 105.000 ;
        RECT 623.725 100.505 624.085 107.065 ;
        RECT 624.865 105.255 625.190 107.120 ;
        RECT 625.505 106.910 625.920 110.260 ;
        RECT 625.530 101.910 625.990 106.595 ;
        RECT 626.315 104.455 626.765 113.275 ;
        RECT 627.175 102.080 627.530 112.385 ;
        RECT 627.840 107.685 628.185 108.740 ;
        RECT 628.500 106.280 628.930 109.270 ;
        RECT 626.245 100.565 626.625 100.945 ;
        RECT 629.135 100.585 629.515 101.960 ;
        RECT 629.905 101.405 630.220 112.455 ;
        RECT 630.920 111.150 631.210 113.210 ;
        RECT 633.705 111.750 634.180 114.800 ;
        RECT 638.660 111.660 639.070 114.755 ;
        RECT 637.700 110.000 638.010 110.030 ;
        RECT 630.840 103.295 631.165 105.665 ;
        RECT 632.490 105.340 632.890 109.305 ;
        RECT 631.575 99.555 631.920 102.015 ;
        RECT 633.210 101.235 633.535 104.000 ;
        RECT 634.195 103.270 634.600 106.600 ;
        RECT 637.700 103.900 638.015 110.000 ;
        RECT 638.845 100.295 639.215 109.395 ;
        RECT 639.790 101.360 640.080 113.195 ;
        RECT 643.240 111.635 643.650 114.730 ;
        RECT 647.695 111.090 648.005 113.605 ;
        RECT 640.685 103.855 641.015 110.050 ;
        RECT 643.605 103.325 644.045 106.600 ;
        RECT 645.985 105.340 646.510 109.280 ;
        RECT 645.145 101.235 645.470 104.000 ;
        RECT 647.660 103.330 648.075 105.720 ;
        RECT 648.690 101.890 649.005 112.575 ;
        RECT 650.020 106.280 650.505 109.290 ;
        RECT 651.200 101.905 651.530 112.600 ;
        RECT 649.390 100.500 649.725 101.850 ;
        RECT 560.980 81.685 561.295 92.735 ;
        RECT 564.815 92.030 565.215 95.080 ;
        RECT 569.735 91.940 570.145 95.035 ;
        RECT 574.315 91.915 574.725 95.010 ;
        RECT 562.650 79.835 562.995 82.295 ;
        RECT 579.765 82.170 580.080 92.855 ;
        RECT 584.950 84.960 585.400 89.120 ;
        RECT 586.650 87.940 587.175 88.380 ;
        RECT 398.050 68.925 398.430 69.305 ;
        RECT 398.040 68.175 398.420 68.555 ;
        RECT 398.085 67.490 398.465 67.870 ;
        RECT 398.050 66.820 398.430 67.200 ;
        RECT 398.765 63.745 399.065 70.785 ;
        RECT 399.885 63.140 400.185 70.070 ;
        RECT 400.540 64.500 400.840 68.560 ;
        RECT 401.195 63.740 401.495 70.090 ;
        RECT 401.790 65.615 402.110 70.775 ;
        RECT 402.510 63.770 402.805 70.595 ;
        RECT 403.640 63.230 403.940 70.040 ;
        RECT 404.430 63.825 404.740 70.015 ;
        RECT 405.225 63.755 405.525 70.585 ;
        RECT 406.350 63.140 406.650 70.080 ;
        RECT 407.030 64.485 407.310 68.575 ;
        RECT 407.800 63.015 408.080 66.050 ;
        RECT 408.560 63.715 408.865 70.075 ;
        RECT 409.410 63.715 409.710 70.535 ;
        RECT 410.550 62.970 410.850 70.125 ;
        RECT 411.215 68.925 411.595 69.305 ;
        RECT 413.485 68.925 413.865 69.330 ;
        RECT 411.220 68.175 411.600 68.555 ;
        RECT 413.490 68.175 413.870 68.580 ;
        RECT 411.220 67.160 411.600 67.540 ;
        RECT 413.005 65.740 413.325 67.870 ;
        RECT 411.435 62.450 411.815 65.470 ;
        RECT 413.615 64.900 413.895 67.305 ;
        RECT 414.225 63.745 414.525 70.785 ;
        RECT 415.345 63.140 415.645 70.070 ;
        RECT 416.000 64.500 416.300 68.560 ;
        RECT 416.655 63.740 416.955 70.090 ;
        RECT 417.250 65.615 417.575 70.775 ;
        RECT 417.970 63.770 418.265 70.595 ;
        RECT 419.100 63.230 419.400 70.040 ;
        RECT 419.890 63.825 420.200 70.015 ;
        RECT 420.685 63.755 420.985 70.585 ;
        RECT 421.810 63.140 422.110 70.080 ;
        RECT 422.490 64.485 422.770 68.575 ;
        RECT 423.260 63.015 423.540 66.050 ;
        RECT 424.020 63.715 424.340 70.075 ;
        RECT 424.870 63.715 425.170 70.535 ;
        RECT 426.010 62.970 426.310 70.125 ;
        RECT 426.950 68.925 427.310 70.755 ;
        RECT 426.645 65.115 427.025 65.495 ;
        RECT 427.350 61.000 427.710 67.560 ;
        RECT 428.490 65.750 428.815 67.615 ;
        RECT 429.130 67.405 429.545 70.755 ;
        RECT 429.155 62.405 429.615 67.090 ;
        RECT 429.940 64.950 430.390 73.770 ;
        RECT 430.800 62.575 431.155 72.880 ;
        RECT 431.465 68.180 431.810 69.235 ;
        RECT 432.125 66.775 432.555 69.765 ;
        RECT 429.870 61.060 430.250 61.440 ;
        RECT 432.760 61.080 433.140 62.455 ;
        RECT 433.530 61.900 433.845 72.950 ;
        RECT 434.545 71.645 434.835 73.705 ;
        RECT 437.330 72.245 437.805 75.295 ;
        RECT 442.285 72.155 442.695 75.250 ;
        RECT 441.325 70.495 441.635 70.525 ;
        RECT 434.465 63.790 434.790 66.160 ;
        RECT 436.115 65.835 436.515 69.800 ;
        RECT 435.200 60.050 435.545 62.510 ;
        RECT 436.835 61.730 437.160 64.495 ;
        RECT 437.820 63.765 438.225 67.095 ;
        RECT 441.325 64.395 441.640 70.495 ;
        RECT 442.470 60.790 442.840 69.890 ;
        RECT 443.415 61.855 443.705 73.690 ;
        RECT 446.865 72.130 447.275 75.225 ;
        RECT 451.320 71.585 451.630 74.100 ;
        RECT 444.310 64.350 444.640 70.545 ;
        RECT 447.230 63.820 447.670 67.095 ;
        RECT 449.610 65.835 450.135 69.775 ;
        RECT 448.770 61.730 449.095 64.495 ;
        RECT 451.285 63.825 451.700 66.215 ;
        RECT 452.315 62.385 452.630 73.070 ;
        RECT 453.645 66.775 454.130 69.785 ;
        RECT 454.825 62.400 455.155 73.095 ;
        RECT 453.015 60.995 453.350 62.345 ;
        RECT 364.660 42.090 364.975 53.140 ;
        RECT 368.495 52.435 368.895 55.485 ;
        RECT 373.415 52.345 373.825 55.440 ;
        RECT 377.995 52.320 378.405 55.415 ;
        RECT 366.330 40.240 366.675 42.700 ;
        RECT 383.445 42.575 383.760 53.260 ;
        RECT 388.630 45.365 389.080 49.525 ;
        RECT 390.330 48.345 390.855 48.785 ;
        RECT 201.570 29.370 201.950 29.750 ;
        RECT 201.560 28.620 201.940 29.000 ;
        RECT 201.605 27.935 201.985 28.315 ;
        RECT 201.570 27.265 201.950 27.645 ;
        RECT 202.285 24.190 202.585 31.230 ;
        RECT 203.405 23.585 203.705 30.515 ;
        RECT 204.060 24.945 204.360 29.005 ;
        RECT 204.715 24.185 205.015 30.535 ;
        RECT 205.310 26.060 205.630 31.220 ;
        RECT 206.030 24.215 206.325 31.040 ;
        RECT 207.160 23.675 207.460 30.485 ;
        RECT 207.950 24.270 208.260 30.460 ;
        RECT 208.745 24.200 209.045 31.030 ;
        RECT 209.870 23.585 210.170 30.525 ;
        RECT 210.550 24.930 210.830 29.020 ;
        RECT 211.320 23.460 211.600 26.495 ;
        RECT 212.080 24.160 212.385 30.520 ;
        RECT 212.930 24.160 213.230 30.980 ;
        RECT 214.070 23.415 214.370 30.570 ;
        RECT 214.735 29.370 215.115 29.750 ;
        RECT 217.005 29.370 217.385 29.775 ;
        RECT 214.740 28.620 215.120 29.000 ;
        RECT 217.010 28.620 217.390 29.025 ;
        RECT 214.740 27.605 215.120 27.985 ;
        RECT 216.525 26.185 216.845 28.315 ;
        RECT 214.955 22.895 215.335 25.915 ;
        RECT 217.135 25.345 217.415 27.750 ;
        RECT 217.745 24.190 218.045 31.230 ;
        RECT 218.865 23.585 219.165 30.515 ;
        RECT 219.520 24.945 219.820 29.005 ;
        RECT 220.175 24.185 220.475 30.535 ;
        RECT 220.770 26.060 221.095 31.220 ;
        RECT 221.490 24.215 221.785 31.040 ;
        RECT 222.620 23.675 222.920 30.485 ;
        RECT 223.410 24.270 223.720 30.460 ;
        RECT 224.205 24.200 224.505 31.030 ;
        RECT 225.330 23.585 225.630 30.525 ;
        RECT 226.010 24.930 226.290 29.020 ;
        RECT 226.780 23.460 227.060 26.495 ;
        RECT 227.540 24.160 227.860 30.520 ;
        RECT 228.390 24.160 228.690 30.980 ;
        RECT 229.530 23.415 229.830 30.570 ;
        RECT 230.470 29.370 230.830 31.200 ;
        RECT 230.165 25.560 230.545 25.940 ;
        RECT 230.870 21.445 231.230 28.005 ;
        RECT 232.010 26.195 232.335 28.060 ;
        RECT 232.650 27.850 233.065 31.200 ;
        RECT 232.675 22.850 233.135 27.535 ;
        RECT 233.460 25.395 233.910 34.215 ;
        RECT 234.320 23.020 234.675 33.325 ;
        RECT 234.985 28.625 235.330 29.680 ;
        RECT 235.645 27.220 236.075 30.210 ;
        RECT 233.390 21.505 233.770 21.885 ;
        RECT 236.280 21.525 236.660 22.900 ;
        RECT 237.050 22.345 237.365 33.395 ;
        RECT 238.065 32.090 238.355 34.150 ;
        RECT 240.850 32.690 241.325 35.740 ;
        RECT 245.805 32.600 246.215 35.695 ;
        RECT 244.845 30.940 245.155 30.970 ;
        RECT 237.985 24.235 238.310 26.605 ;
        RECT 239.635 26.280 240.035 30.245 ;
        RECT 238.720 20.495 239.065 22.955 ;
        RECT 240.355 22.175 240.680 24.940 ;
        RECT 241.340 24.210 241.745 27.540 ;
        RECT 244.845 24.840 245.160 30.940 ;
        RECT 245.990 21.235 246.360 30.335 ;
        RECT 246.935 22.300 247.225 34.135 ;
        RECT 250.385 32.575 250.795 35.670 ;
        RECT 254.840 32.030 255.150 34.545 ;
        RECT 247.830 24.795 248.160 30.990 ;
        RECT 250.750 24.265 251.190 27.540 ;
        RECT 253.130 26.280 253.655 30.220 ;
        RECT 252.290 22.175 252.615 24.940 ;
        RECT 254.805 24.270 255.220 26.660 ;
        RECT 255.835 22.830 256.150 33.515 ;
        RECT 257.165 27.220 257.650 30.230 ;
        RECT 258.345 22.845 258.675 33.540 ;
        RECT 263.625 29.140 266.950 29.730 ;
        RECT 263.625 28.525 264.375 29.140 ;
        RECT 265.530 25.685 266.200 28.335 ;
        RECT 256.535 21.440 256.870 22.790 ;
        RECT 267.490 9.530 267.940 28.570 ;
        RECT 269.280 8.755 269.695 29.935 ;
        RECT 273.020 22.355 273.375 33.440 ;
        RECT 276.765 32.080 277.055 34.140 ;
        RECT 279.535 32.680 280.035 35.730 ;
        RECT 284.505 32.590 284.915 35.685 ;
        RECT 283.545 30.930 283.855 30.960 ;
        RECT 274.345 27.210 274.815 30.200 ;
        RECT 276.695 24.225 277.010 26.595 ;
        RECT 278.315 26.270 278.735 30.235 ;
        RECT 274.980 21.515 275.360 22.890 ;
        RECT 277.420 20.485 277.765 22.945 ;
        RECT 279.055 22.165 279.380 24.930 ;
        RECT 280.040 24.200 280.445 27.530 ;
        RECT 283.545 24.830 283.860 30.930 ;
        RECT 284.690 21.225 285.060 30.325 ;
        RECT 285.635 22.290 285.925 34.125 ;
        RECT 289.085 32.565 289.495 35.660 ;
        RECT 293.540 32.020 293.850 34.535 ;
        RECT 297.790 33.720 298.170 34.100 ;
        RECT 299.920 33.720 300.300 34.100 ;
        RECT 286.530 24.785 286.860 30.980 ;
        RECT 289.435 24.255 289.890 27.530 ;
        RECT 291.795 26.270 292.340 30.210 ;
        RECT 295.850 27.210 296.285 30.220 ;
        RECT 290.990 22.165 291.315 24.930 ;
        RECT 293.505 24.260 293.920 26.650 ;
        RECT 297.045 22.835 297.375 33.530 ;
        RECT 298.480 27.170 298.865 32.955 ;
        RECT 295.235 21.430 295.570 22.780 ;
        RECT 298.840 22.415 299.265 26.690 ;
        RECT 300.540 24.180 300.840 31.220 ;
        RECT 301.660 23.575 301.960 30.505 ;
        RECT 302.970 24.175 303.270 30.525 ;
        RECT 297.500 21.505 297.880 21.885 ;
        RECT 299.695 21.490 300.075 21.870 ;
        RECT 303.565 21.430 303.855 31.210 ;
        RECT 304.285 24.205 304.580 31.030 ;
        RECT 305.415 23.665 305.715 30.475 ;
        RECT 306.205 24.260 306.515 34.300 ;
        RECT 315.395 32.545 315.775 32.925 ;
        RECT 307.000 24.190 307.300 31.020 ;
        RECT 308.125 23.575 308.425 30.515 ;
        RECT 309.575 23.450 309.855 26.485 ;
        RECT 310.335 24.150 310.615 30.510 ;
        RECT 311.185 24.150 311.485 30.970 ;
        RECT 312.325 23.405 312.625 30.560 ;
        RECT 312.970 27.595 313.350 27.975 ;
        RECT 312.970 25.540 313.350 25.920 ;
        RECT 314.820 25.420 315.135 29.745 ;
        RECT 315.430 27.495 315.710 29.025 ;
        RECT 316.000 24.180 316.300 31.220 ;
        RECT 317.120 23.575 317.420 30.505 ;
        RECT 317.775 24.935 318.075 28.995 ;
        RECT 318.430 24.175 318.730 30.525 ;
        RECT 315.295 22.370 315.675 22.750 ;
        RECT 319.025 21.965 319.315 31.210 ;
        RECT 319.745 24.205 320.040 31.030 ;
        RECT 320.875 23.665 321.175 30.475 ;
        RECT 321.665 24.260 321.975 32.995 ;
        RECT 322.460 24.190 322.760 31.020 ;
        RECT 323.585 23.575 323.885 30.515 ;
        RECT 324.265 24.920 324.545 29.010 ;
        RECT 325.035 23.450 325.315 26.485 ;
        RECT 325.795 24.150 326.075 30.510 ;
        RECT 326.645 24.150 326.945 30.970 ;
        RECT 327.785 23.405 328.085 30.560 ;
        RECT 329.710 29.325 330.085 37.165 ;
        RECT 331.565 28.575 331.865 39.115 ;
        RECT 332.880 27.395 333.260 37.650 ;
        RECT 333.750 25.240 334.185 38.815 ;
        RECT 389.460 38.080 389.975 48.130 ;
        RECT 391.145 36.725 391.730 47.505 ;
        RECT 392.735 45.025 393.090 58.935 ;
        RECT 456.080 58.305 456.530 68.570 ;
        RECT 394.360 45.945 394.720 57.335 ;
        RECT 457.245 56.765 457.730 65.650 ;
        RECT 464.075 56.120 464.480 68.000 ;
        RECT 466.150 58.020 466.540 69.600 ;
        RECT 469.420 61.940 469.775 73.025 ;
        RECT 473.165 71.665 473.455 73.725 ;
        RECT 475.935 72.265 476.435 75.315 ;
        RECT 480.905 72.175 481.315 75.270 ;
        RECT 479.945 70.515 480.255 70.545 ;
        RECT 470.745 66.795 471.215 69.785 ;
        RECT 473.095 63.810 473.410 66.180 ;
        RECT 474.715 65.855 475.135 69.820 ;
        RECT 471.380 61.100 471.760 62.475 ;
        RECT 473.820 60.070 474.165 62.530 ;
        RECT 475.455 61.750 475.780 64.515 ;
        RECT 476.440 63.785 476.845 67.115 ;
        RECT 479.945 64.415 480.260 70.515 ;
        RECT 481.090 60.810 481.460 69.910 ;
        RECT 482.035 61.875 482.325 73.710 ;
        RECT 485.485 72.150 485.895 75.245 ;
        RECT 489.940 71.605 490.250 74.120 ;
        RECT 494.190 73.305 494.570 73.685 ;
        RECT 496.320 73.305 496.700 73.685 ;
        RECT 482.930 64.370 483.260 70.565 ;
        RECT 485.835 63.840 486.290 67.115 ;
        RECT 488.195 65.855 488.740 69.795 ;
        RECT 492.250 66.795 492.685 69.805 ;
        RECT 487.390 61.750 487.715 64.515 ;
        RECT 489.905 63.845 490.320 66.235 ;
        RECT 493.445 62.420 493.775 73.115 ;
        RECT 494.880 66.755 495.265 72.540 ;
        RECT 491.635 61.015 491.970 62.365 ;
        RECT 495.240 62.000 495.665 66.275 ;
        RECT 496.940 63.765 497.240 70.805 ;
        RECT 498.060 63.160 498.360 70.090 ;
        RECT 499.370 63.760 499.670 70.110 ;
        RECT 493.900 61.090 494.280 61.470 ;
        RECT 496.095 61.075 496.475 61.455 ;
        RECT 499.965 61.015 500.255 70.795 ;
        RECT 500.685 63.790 500.980 70.615 ;
        RECT 501.815 63.250 502.115 70.060 ;
        RECT 502.605 63.845 502.915 73.885 ;
        RECT 511.795 72.130 512.175 72.510 ;
        RECT 503.400 63.775 503.700 70.605 ;
        RECT 504.525 63.160 504.825 70.100 ;
        RECT 505.975 63.035 506.255 66.070 ;
        RECT 506.735 63.735 507.015 70.095 ;
        RECT 507.585 63.735 507.885 70.555 ;
        RECT 508.725 62.990 509.025 70.145 ;
        RECT 509.370 67.180 509.750 67.560 ;
        RECT 509.370 65.125 509.750 65.505 ;
        RECT 511.220 65.005 511.535 69.330 ;
        RECT 511.830 67.080 512.110 68.610 ;
        RECT 512.400 63.765 512.700 70.805 ;
        RECT 513.520 63.160 513.820 70.090 ;
        RECT 514.175 64.520 514.475 68.580 ;
        RECT 514.830 63.760 515.130 70.110 ;
        RECT 511.695 61.955 512.075 62.335 ;
        RECT 515.425 61.550 515.715 70.795 ;
        RECT 516.145 63.790 516.440 70.615 ;
        RECT 517.275 63.250 517.575 70.060 ;
        RECT 518.065 63.845 518.375 72.580 ;
        RECT 518.860 63.775 519.160 70.605 ;
        RECT 519.985 63.160 520.285 70.100 ;
        RECT 520.665 64.505 520.945 68.595 ;
        RECT 521.435 63.035 521.715 66.070 ;
        RECT 522.195 63.735 522.475 70.095 ;
        RECT 523.045 63.735 523.345 70.555 ;
        RECT 524.185 62.990 524.485 70.145 ;
        RECT 526.265 68.865 526.640 77.145 ;
        RECT 528.010 68.025 528.310 79.135 ;
        RECT 529.200 67.075 529.580 77.330 ;
        RECT 530.070 64.920 530.505 78.495 ;
        RECT 585.780 77.695 586.295 87.745 ;
        RECT 587.465 76.340 588.050 87.120 ;
        RECT 589.320 84.585 589.675 98.375 ;
        RECT 652.665 97.745 653.115 108.235 ;
        RECT 590.945 85.490 591.305 96.775 ;
        RECT 653.830 96.205 654.315 105.365 ;
        RECT 660.290 96.015 660.695 107.545 ;
        RECT 662.365 97.915 662.755 109.015 ;
        RECT 665.770 101.445 666.125 112.530 ;
        RECT 669.515 111.170 669.805 113.230 ;
        RECT 672.285 111.770 672.785 114.820 ;
        RECT 677.255 111.680 677.665 114.775 ;
        RECT 676.295 110.020 676.605 110.050 ;
        RECT 667.095 106.300 667.565 109.290 ;
        RECT 669.445 103.315 669.760 105.685 ;
        RECT 671.065 105.360 671.485 109.325 ;
        RECT 667.730 100.605 668.110 101.980 ;
        RECT 670.170 99.575 670.515 102.035 ;
        RECT 671.805 101.255 672.130 104.020 ;
        RECT 672.790 103.290 673.195 106.620 ;
        RECT 676.295 103.920 676.610 110.020 ;
        RECT 677.440 100.315 677.810 109.415 ;
        RECT 678.385 101.380 678.675 113.215 ;
        RECT 681.835 111.655 682.245 114.750 ;
        RECT 686.290 111.110 686.600 113.625 ;
        RECT 690.540 112.810 690.920 113.190 ;
        RECT 692.670 112.810 693.050 113.190 ;
        RECT 679.280 103.875 679.610 110.070 ;
        RECT 682.185 103.345 682.640 106.620 ;
        RECT 684.545 105.360 685.090 109.300 ;
        RECT 688.600 106.300 689.035 109.310 ;
        RECT 683.740 101.255 684.065 104.020 ;
        RECT 686.255 103.350 686.670 105.740 ;
        RECT 689.795 101.925 690.125 112.620 ;
        RECT 691.230 106.260 691.615 112.045 ;
        RECT 687.985 100.520 688.320 101.870 ;
        RECT 691.590 101.505 692.015 105.780 ;
        RECT 693.290 103.270 693.590 110.310 ;
        RECT 694.410 102.665 694.710 109.595 ;
        RECT 695.720 103.265 696.020 109.615 ;
        RECT 690.250 100.595 690.630 100.975 ;
        RECT 692.445 100.580 692.825 100.960 ;
        RECT 696.315 100.520 696.605 110.300 ;
        RECT 697.035 103.295 697.330 110.120 ;
        RECT 698.165 102.755 698.465 109.565 ;
        RECT 698.955 103.350 699.265 113.390 ;
        RECT 708.145 111.635 708.525 112.015 ;
        RECT 699.750 103.280 700.050 110.110 ;
        RECT 700.875 102.665 701.175 109.605 ;
        RECT 702.325 102.540 702.605 105.575 ;
        RECT 703.085 103.240 703.365 109.600 ;
        RECT 703.935 103.240 704.235 110.060 ;
        RECT 705.075 102.495 705.375 109.650 ;
        RECT 705.720 106.685 706.100 107.065 ;
        RECT 705.720 104.630 706.100 105.010 ;
        RECT 707.570 104.510 707.885 108.835 ;
        RECT 708.180 106.585 708.460 108.115 ;
        RECT 708.750 103.270 709.050 110.310 ;
        RECT 709.870 102.665 710.170 109.595 ;
        RECT 710.525 104.025 710.825 108.085 ;
        RECT 711.180 103.265 711.480 109.615 ;
        RECT 708.045 101.460 708.425 101.840 ;
        RECT 711.775 101.055 712.065 110.300 ;
        RECT 712.495 103.295 712.790 110.120 ;
        RECT 713.625 102.755 713.925 109.565 ;
        RECT 714.415 103.350 714.725 112.085 ;
        RECT 715.210 103.280 715.510 110.110 ;
        RECT 716.335 102.665 716.635 109.605 ;
        RECT 717.015 104.010 717.295 108.100 ;
        RECT 717.785 102.540 718.065 105.575 ;
        RECT 718.545 103.240 718.825 109.600 ;
        RECT 719.395 103.240 719.695 110.060 ;
        RECT 720.535 102.495 720.835 109.650 ;
        RECT 722.740 108.420 723.115 116.620 ;
        RECT 724.485 107.615 724.785 118.610 ;
        RECT 725.565 106.545 725.945 116.800 ;
        RECT 726.435 104.390 726.870 117.965 ;
        RECT 782.290 117.245 782.805 127.295 ;
        RECT 783.975 115.890 784.560 126.670 ;
        RECT 785.495 124.150 785.850 138.205 ;
        RECT 848.840 137.575 849.290 147.690 ;
        RECT 787.120 124.955 787.480 136.605 ;
        RECT 850.005 136.035 850.490 144.790 ;
        RECT 856.610 135.410 857.015 146.940 ;
        RECT 858.685 137.310 859.075 148.410 ;
        RECT 861.955 140.885 862.310 151.970 ;
        RECT 865.700 150.610 865.990 152.670 ;
        RECT 868.470 151.210 868.970 154.260 ;
        RECT 873.440 151.120 873.850 154.215 ;
        RECT 872.480 149.460 872.790 149.490 ;
        RECT 863.280 145.740 863.750 148.730 ;
        RECT 865.630 142.755 865.945 145.125 ;
        RECT 867.250 144.800 867.670 148.765 ;
        RECT 863.915 140.045 864.295 141.420 ;
        RECT 866.355 139.015 866.700 141.475 ;
        RECT 867.990 140.695 868.315 143.460 ;
        RECT 868.975 142.730 869.380 146.060 ;
        RECT 872.480 143.360 872.795 149.460 ;
        RECT 873.625 139.755 873.995 148.855 ;
        RECT 874.570 140.820 874.860 152.655 ;
        RECT 878.020 151.095 878.430 154.190 ;
        RECT 882.475 150.550 882.785 153.065 ;
        RECT 886.725 152.250 887.105 152.630 ;
        RECT 888.855 152.250 889.235 152.630 ;
        RECT 875.465 143.315 875.795 149.510 ;
        RECT 878.370 142.785 878.825 146.060 ;
        RECT 880.730 144.800 881.275 148.740 ;
        RECT 884.785 145.740 885.220 148.750 ;
        RECT 879.925 140.695 880.250 143.460 ;
        RECT 882.440 142.790 882.855 145.180 ;
        RECT 885.980 141.365 886.310 152.060 ;
        RECT 887.415 145.700 887.800 151.485 ;
        RECT 884.170 139.960 884.505 141.310 ;
        RECT 887.775 140.945 888.200 145.220 ;
        RECT 889.475 142.710 889.775 149.750 ;
        RECT 890.595 142.105 890.895 149.035 ;
        RECT 891.905 142.705 892.205 149.055 ;
        RECT 886.435 140.035 886.815 140.415 ;
        RECT 888.630 140.020 889.010 140.400 ;
        RECT 892.500 139.960 892.790 149.740 ;
        RECT 893.220 142.735 893.515 149.560 ;
        RECT 894.350 142.195 894.650 149.005 ;
        RECT 895.140 142.790 895.450 152.830 ;
        RECT 904.330 151.075 904.710 151.455 ;
        RECT 895.935 142.720 896.235 149.550 ;
        RECT 897.060 142.105 897.360 149.045 ;
        RECT 898.510 141.980 898.790 145.015 ;
        RECT 899.270 142.680 899.550 149.040 ;
        RECT 900.120 142.680 900.420 149.500 ;
        RECT 901.260 141.935 901.560 149.090 ;
        RECT 901.905 146.125 902.285 146.505 ;
        RECT 901.905 144.070 902.285 144.450 ;
        RECT 903.755 143.950 904.070 148.275 ;
        RECT 904.365 146.025 904.645 147.555 ;
        RECT 904.935 142.710 905.235 149.750 ;
        RECT 906.055 142.105 906.355 149.035 ;
        RECT 906.710 143.465 907.010 147.525 ;
        RECT 907.365 142.705 907.665 149.055 ;
        RECT 904.230 140.900 904.610 141.280 ;
        RECT 907.960 140.495 908.250 149.740 ;
        RECT 908.680 142.735 908.975 149.560 ;
        RECT 909.810 142.195 910.110 149.005 ;
        RECT 910.600 142.790 910.910 151.525 ;
        RECT 911.395 142.720 911.695 149.550 ;
        RECT 912.520 142.105 912.820 149.045 ;
        RECT 913.200 143.450 913.480 147.540 ;
        RECT 913.970 141.980 914.250 145.015 ;
        RECT 914.730 142.680 915.010 149.040 ;
        RECT 915.580 142.680 915.880 149.500 ;
        RECT 916.720 141.935 917.020 149.090 ;
        RECT 918.760 147.830 919.135 156.030 ;
        RECT 920.505 147.025 920.805 158.020 ;
        RECT 921.950 145.970 922.330 156.225 ;
        RECT 922.820 143.815 923.255 157.390 ;
        RECT 978.525 156.635 979.040 166.685 ;
        RECT 987.190 166.235 987.570 166.615 ;
        RECT 980.210 155.280 980.795 166.060 ;
        RECT 987.155 165.565 987.535 165.945 ;
        RECT 987.870 162.490 988.170 169.530 ;
        RECT 988.990 161.885 989.290 168.815 ;
        RECT 989.645 163.245 989.945 167.305 ;
        RECT 990.300 162.485 990.600 168.835 ;
        RECT 990.895 164.360 991.215 169.520 ;
        RECT 991.615 162.515 991.910 169.340 ;
        RECT 992.745 161.975 993.045 168.785 ;
        RECT 993.535 162.570 993.845 168.760 ;
        RECT 994.330 162.500 994.630 169.330 ;
        RECT 995.455 161.885 995.755 168.825 ;
        RECT 996.135 163.230 996.415 167.320 ;
        RECT 996.905 161.760 997.185 164.795 ;
        RECT 997.665 162.460 997.970 168.820 ;
        RECT 998.515 162.460 998.815 169.280 ;
        RECT 999.655 161.715 999.955 168.870 ;
        RECT 1000.320 167.670 1000.700 168.050 ;
        RECT 1002.590 167.670 1002.970 168.075 ;
        RECT 1000.325 166.920 1000.705 167.300 ;
        RECT 1002.595 166.920 1002.975 167.325 ;
        RECT 1000.325 165.905 1000.705 166.285 ;
        RECT 1002.110 164.485 1002.430 166.615 ;
        RECT 1000.540 161.195 1000.920 164.215 ;
        RECT 1002.720 163.645 1003.000 166.050 ;
        RECT 1003.330 162.490 1003.630 169.530 ;
        RECT 1004.450 161.885 1004.750 168.815 ;
        RECT 1005.105 163.245 1005.405 167.305 ;
        RECT 1005.760 162.485 1006.060 168.835 ;
        RECT 1006.355 164.360 1006.680 169.520 ;
        RECT 1007.075 162.515 1007.370 169.340 ;
        RECT 1008.205 161.975 1008.505 168.785 ;
        RECT 1008.995 162.570 1009.305 168.760 ;
        RECT 1009.790 162.500 1010.090 169.330 ;
        RECT 1010.915 161.885 1011.215 168.825 ;
        RECT 1011.595 163.230 1011.875 167.320 ;
        RECT 1012.365 161.760 1012.645 164.795 ;
        RECT 1013.125 162.460 1013.445 168.820 ;
        RECT 1013.975 162.460 1014.275 169.280 ;
        RECT 1015.115 161.715 1015.415 168.870 ;
        RECT 1016.055 167.670 1016.415 169.500 ;
        RECT 1015.750 163.860 1016.130 164.240 ;
        RECT 1016.455 159.745 1016.815 166.305 ;
        RECT 1017.595 164.495 1017.920 166.360 ;
        RECT 1018.235 166.150 1018.650 169.500 ;
        RECT 1018.260 161.150 1018.720 165.835 ;
        RECT 1019.045 163.695 1019.495 172.515 ;
        RECT 1019.905 161.320 1020.260 171.625 ;
        RECT 1020.570 166.925 1020.915 167.980 ;
        RECT 1021.230 165.520 1021.660 168.510 ;
        RECT 1018.975 159.805 1019.355 160.185 ;
        RECT 1021.865 159.825 1022.245 161.200 ;
        RECT 1022.635 160.645 1022.950 171.695 ;
        RECT 1023.650 170.390 1023.940 172.450 ;
        RECT 1026.435 170.990 1026.910 174.040 ;
        RECT 1031.390 170.900 1031.800 173.995 ;
        RECT 1030.430 169.240 1030.740 169.270 ;
        RECT 1023.570 162.535 1023.895 164.905 ;
        RECT 1025.220 164.580 1025.620 168.545 ;
        RECT 1024.305 158.795 1024.650 161.255 ;
        RECT 1025.940 160.475 1026.265 163.240 ;
        RECT 1026.925 162.510 1027.330 165.840 ;
        RECT 1030.430 163.140 1030.745 169.240 ;
        RECT 1031.575 159.535 1031.945 168.635 ;
        RECT 1032.520 160.600 1032.810 172.435 ;
        RECT 1035.970 170.875 1036.380 173.970 ;
        RECT 1040.425 170.330 1040.735 172.845 ;
        RECT 1033.415 163.095 1033.745 169.290 ;
        RECT 1036.335 162.565 1036.775 165.840 ;
        RECT 1038.715 164.580 1039.240 168.520 ;
        RECT 1037.875 160.475 1038.200 163.240 ;
        RECT 1040.390 162.570 1040.805 164.960 ;
        RECT 1041.420 161.130 1041.735 171.815 ;
        RECT 1042.750 165.520 1043.235 168.530 ;
        RECT 1043.930 161.145 1044.260 171.840 ;
        RECT 1042.120 159.740 1042.455 161.090 ;
        RECT 953.710 140.975 954.025 152.025 ;
        RECT 957.545 151.320 957.945 154.370 ;
        RECT 962.465 151.230 962.875 154.325 ;
        RECT 967.045 151.205 967.455 154.300 ;
        RECT 955.380 139.125 955.725 141.585 ;
        RECT 972.495 141.460 972.810 152.145 ;
        RECT 977.680 144.250 978.130 148.410 ;
        RECT 979.380 147.230 979.905 147.670 ;
        RECT 790.960 128.270 791.340 128.650 ;
        RECT 790.950 127.520 791.330 127.900 ;
        RECT 790.995 126.835 791.375 127.215 ;
        RECT 790.960 126.165 791.340 126.545 ;
        RECT 791.675 123.090 791.975 130.130 ;
        RECT 792.795 122.485 793.095 129.415 ;
        RECT 793.450 123.845 793.750 127.905 ;
        RECT 794.105 123.085 794.405 129.435 ;
        RECT 794.700 124.960 795.020 130.120 ;
        RECT 795.420 123.115 795.715 129.940 ;
        RECT 796.550 122.575 796.850 129.385 ;
        RECT 797.340 123.170 797.650 129.360 ;
        RECT 798.135 123.100 798.435 129.930 ;
        RECT 799.260 122.485 799.560 129.425 ;
        RECT 799.940 123.830 800.220 127.920 ;
        RECT 800.710 122.360 800.990 125.395 ;
        RECT 801.470 123.060 801.775 129.420 ;
        RECT 802.320 123.060 802.620 129.880 ;
        RECT 803.460 122.315 803.760 129.470 ;
        RECT 804.125 128.270 804.505 128.650 ;
        RECT 806.395 128.270 806.775 128.675 ;
        RECT 804.130 127.520 804.510 127.900 ;
        RECT 806.400 127.520 806.780 127.925 ;
        RECT 804.130 126.505 804.510 126.885 ;
        RECT 805.915 125.085 806.235 127.215 ;
        RECT 804.345 121.795 804.725 124.815 ;
        RECT 806.525 124.245 806.805 126.650 ;
        RECT 807.135 123.090 807.435 130.130 ;
        RECT 808.255 122.485 808.555 129.415 ;
        RECT 808.910 123.845 809.210 127.905 ;
        RECT 809.565 123.085 809.865 129.435 ;
        RECT 810.160 124.960 810.485 130.120 ;
        RECT 810.880 123.115 811.175 129.940 ;
        RECT 812.010 122.575 812.310 129.385 ;
        RECT 812.800 123.170 813.110 129.360 ;
        RECT 813.595 123.100 813.895 129.930 ;
        RECT 814.720 122.485 815.020 129.425 ;
        RECT 815.400 123.830 815.680 127.920 ;
        RECT 816.170 122.360 816.450 125.395 ;
        RECT 816.930 123.060 817.250 129.420 ;
        RECT 817.780 123.060 818.080 129.880 ;
        RECT 818.920 122.315 819.220 129.470 ;
        RECT 819.860 128.270 820.220 130.100 ;
        RECT 819.555 124.460 819.935 124.840 ;
        RECT 820.260 120.345 820.620 126.905 ;
        RECT 821.400 125.095 821.725 126.960 ;
        RECT 822.040 126.750 822.455 130.100 ;
        RECT 822.065 121.750 822.525 126.435 ;
        RECT 822.850 124.295 823.300 133.115 ;
        RECT 823.710 121.920 824.065 132.225 ;
        RECT 824.375 127.525 824.720 128.580 ;
        RECT 825.035 126.120 825.465 129.110 ;
        RECT 822.780 120.405 823.160 120.785 ;
        RECT 825.670 120.425 826.050 121.800 ;
        RECT 826.440 121.245 826.755 132.295 ;
        RECT 827.455 130.990 827.745 133.050 ;
        RECT 830.240 131.590 830.715 134.640 ;
        RECT 835.195 131.500 835.605 134.595 ;
        RECT 834.235 129.840 834.545 129.870 ;
        RECT 827.375 123.135 827.700 125.505 ;
        RECT 829.025 125.180 829.425 129.145 ;
        RECT 828.110 119.395 828.455 121.855 ;
        RECT 829.745 121.075 830.070 123.840 ;
        RECT 830.730 123.110 831.135 126.440 ;
        RECT 834.235 123.740 834.550 129.840 ;
        RECT 835.380 120.135 835.750 129.235 ;
        RECT 836.325 121.200 836.615 133.035 ;
        RECT 839.775 131.475 840.185 134.570 ;
        RECT 844.230 130.930 844.540 133.445 ;
        RECT 837.220 123.695 837.550 129.890 ;
        RECT 840.140 123.165 840.580 126.440 ;
        RECT 842.520 125.180 843.045 129.120 ;
        RECT 841.680 121.075 842.005 123.840 ;
        RECT 844.195 123.170 844.610 125.560 ;
        RECT 845.225 121.730 845.540 132.415 ;
        RECT 846.555 126.120 847.040 129.130 ;
        RECT 847.735 121.745 848.065 132.440 ;
        RECT 845.925 120.340 846.260 121.690 ;
        RECT 757.315 101.415 757.630 112.465 ;
        RECT 761.150 111.760 761.550 114.810 ;
        RECT 766.070 111.670 766.480 114.765 ;
        RECT 770.650 111.645 771.060 114.740 ;
        RECT 758.985 99.565 759.330 102.025 ;
        RECT 776.100 101.900 776.415 112.585 ;
        RECT 781.285 104.690 781.735 108.850 ;
        RECT 782.985 107.670 783.510 108.110 ;
        RECT 594.295 88.720 594.675 89.100 ;
        RECT 594.285 87.970 594.665 88.350 ;
        RECT 594.330 87.285 594.710 87.665 ;
        RECT 594.295 86.615 594.675 86.995 ;
        RECT 595.010 83.540 595.310 90.580 ;
        RECT 596.130 82.935 596.430 89.865 ;
        RECT 596.785 84.295 597.085 88.355 ;
        RECT 597.440 83.535 597.740 89.885 ;
        RECT 598.035 85.410 598.355 90.570 ;
        RECT 598.755 83.565 599.050 90.390 ;
        RECT 599.885 83.025 600.185 89.835 ;
        RECT 600.675 83.620 600.985 89.810 ;
        RECT 601.470 83.550 601.770 90.380 ;
        RECT 602.595 82.935 602.895 89.875 ;
        RECT 603.275 84.280 603.555 88.370 ;
        RECT 604.045 82.810 604.325 85.845 ;
        RECT 604.805 83.510 605.110 89.870 ;
        RECT 605.655 83.510 605.955 90.330 ;
        RECT 606.795 82.765 607.095 89.920 ;
        RECT 607.460 88.720 607.840 89.100 ;
        RECT 609.730 88.720 610.110 89.125 ;
        RECT 607.465 87.970 607.845 88.350 ;
        RECT 609.735 87.970 610.115 88.375 ;
        RECT 607.465 86.955 607.845 87.335 ;
        RECT 609.250 85.535 609.570 87.665 ;
        RECT 607.680 82.245 608.060 85.265 ;
        RECT 609.860 84.695 610.140 87.100 ;
        RECT 610.470 83.540 610.770 90.580 ;
        RECT 611.590 82.935 611.890 89.865 ;
        RECT 612.245 84.295 612.545 88.355 ;
        RECT 612.900 83.535 613.200 89.885 ;
        RECT 613.495 85.410 613.820 90.570 ;
        RECT 614.215 83.565 614.510 90.390 ;
        RECT 615.345 83.025 615.645 89.835 ;
        RECT 616.135 83.620 616.445 89.810 ;
        RECT 616.930 83.550 617.230 90.380 ;
        RECT 618.055 82.935 618.355 89.875 ;
        RECT 618.735 84.280 619.015 88.370 ;
        RECT 619.505 82.810 619.785 85.845 ;
        RECT 620.265 83.510 620.585 89.870 ;
        RECT 621.115 83.510 621.415 90.330 ;
        RECT 622.255 82.765 622.555 89.920 ;
        RECT 623.195 88.720 623.555 90.550 ;
        RECT 622.890 84.910 623.270 85.290 ;
        RECT 623.595 80.795 623.955 87.355 ;
        RECT 624.735 85.545 625.060 87.410 ;
        RECT 625.375 87.200 625.790 90.550 ;
        RECT 625.400 82.200 625.860 86.885 ;
        RECT 626.185 84.745 626.635 93.565 ;
        RECT 627.045 82.370 627.400 92.675 ;
        RECT 627.710 87.975 628.055 89.030 ;
        RECT 628.370 86.570 628.800 89.560 ;
        RECT 626.115 80.855 626.495 81.235 ;
        RECT 629.005 80.875 629.385 82.250 ;
        RECT 629.775 81.695 630.090 92.745 ;
        RECT 630.790 91.440 631.080 93.500 ;
        RECT 633.575 92.040 634.050 95.090 ;
        RECT 638.530 91.950 638.940 95.045 ;
        RECT 637.570 90.290 637.880 90.320 ;
        RECT 630.710 83.585 631.035 85.955 ;
        RECT 632.360 85.630 632.760 89.595 ;
        RECT 631.445 79.845 631.790 82.305 ;
        RECT 633.080 81.525 633.405 84.290 ;
        RECT 634.065 83.560 634.470 86.890 ;
        RECT 637.570 84.190 637.885 90.290 ;
        RECT 638.715 80.585 639.085 89.685 ;
        RECT 639.660 81.650 639.950 93.485 ;
        RECT 643.110 91.925 643.520 95.020 ;
        RECT 647.565 91.380 647.875 93.895 ;
        RECT 640.555 84.145 640.885 90.340 ;
        RECT 643.475 83.615 643.915 86.890 ;
        RECT 645.855 85.630 646.380 89.570 ;
        RECT 645.015 81.525 645.340 84.290 ;
        RECT 647.530 83.620 647.945 86.010 ;
        RECT 648.560 82.180 648.875 92.865 ;
        RECT 649.890 86.570 650.375 89.580 ;
        RECT 651.070 82.195 651.400 92.890 ;
        RECT 649.260 80.790 649.595 82.140 ;
        RECT 560.910 61.855 561.225 72.905 ;
        RECT 564.745 72.200 565.145 75.250 ;
        RECT 569.665 72.110 570.075 75.205 ;
        RECT 574.245 72.085 574.655 75.180 ;
        RECT 562.580 60.005 562.925 62.465 ;
        RECT 579.695 62.340 580.010 73.025 ;
        RECT 584.880 65.130 585.330 69.290 ;
        RECT 586.580 68.110 587.105 68.550 ;
        RECT 398.000 49.115 398.380 49.495 ;
        RECT 397.990 48.365 398.370 48.745 ;
        RECT 398.035 47.680 398.415 48.060 ;
        RECT 398.000 47.010 398.380 47.390 ;
        RECT 398.715 43.935 399.015 50.975 ;
        RECT 399.835 43.330 400.135 50.260 ;
        RECT 400.490 44.690 400.790 48.750 ;
        RECT 401.145 43.930 401.445 50.280 ;
        RECT 401.740 45.805 402.060 50.965 ;
        RECT 402.460 43.960 402.755 50.785 ;
        RECT 403.590 43.420 403.890 50.230 ;
        RECT 404.380 44.015 404.690 50.205 ;
        RECT 405.175 43.945 405.475 50.775 ;
        RECT 406.300 43.330 406.600 50.270 ;
        RECT 406.980 44.675 407.260 48.765 ;
        RECT 407.750 43.205 408.030 46.240 ;
        RECT 408.510 43.905 408.815 50.265 ;
        RECT 409.360 43.905 409.660 50.725 ;
        RECT 410.500 43.160 410.800 50.315 ;
        RECT 411.165 49.115 411.545 49.495 ;
        RECT 413.435 49.115 413.815 49.520 ;
        RECT 411.170 48.365 411.550 48.745 ;
        RECT 413.440 48.365 413.820 48.770 ;
        RECT 411.170 47.350 411.550 47.730 ;
        RECT 412.955 45.930 413.275 48.060 ;
        RECT 411.385 42.640 411.765 45.660 ;
        RECT 413.565 45.090 413.845 47.495 ;
        RECT 414.175 43.935 414.475 50.975 ;
        RECT 415.295 43.330 415.595 50.260 ;
        RECT 415.950 44.690 416.250 48.750 ;
        RECT 416.605 43.930 416.905 50.280 ;
        RECT 417.200 45.805 417.525 50.965 ;
        RECT 417.920 43.960 418.215 50.785 ;
        RECT 419.050 43.420 419.350 50.230 ;
        RECT 419.840 44.015 420.150 50.205 ;
        RECT 420.635 43.945 420.935 50.775 ;
        RECT 421.760 43.330 422.060 50.270 ;
        RECT 422.440 44.675 422.720 48.765 ;
        RECT 423.210 43.205 423.490 46.240 ;
        RECT 423.970 43.905 424.290 50.265 ;
        RECT 424.820 43.905 425.120 50.725 ;
        RECT 425.960 43.160 426.260 50.315 ;
        RECT 426.900 49.115 427.260 50.945 ;
        RECT 426.595 45.305 426.975 45.685 ;
        RECT 427.300 41.190 427.660 47.750 ;
        RECT 428.440 45.940 428.765 47.805 ;
        RECT 429.080 47.595 429.495 50.945 ;
        RECT 429.105 42.595 429.565 47.280 ;
        RECT 429.890 45.140 430.340 53.960 ;
        RECT 430.750 42.765 431.105 53.070 ;
        RECT 431.415 48.370 431.760 49.425 ;
        RECT 432.075 46.965 432.505 49.955 ;
        RECT 429.820 41.250 430.200 41.630 ;
        RECT 432.710 41.270 433.090 42.645 ;
        RECT 433.480 42.090 433.795 53.140 ;
        RECT 434.495 51.835 434.785 53.895 ;
        RECT 437.280 52.435 437.755 55.485 ;
        RECT 442.235 52.345 442.645 55.440 ;
        RECT 441.275 50.685 441.585 50.715 ;
        RECT 434.415 43.980 434.740 46.350 ;
        RECT 436.065 46.025 436.465 49.990 ;
        RECT 435.150 40.240 435.495 42.700 ;
        RECT 436.785 41.920 437.110 44.685 ;
        RECT 437.770 43.955 438.175 47.285 ;
        RECT 441.275 44.585 441.590 50.685 ;
        RECT 442.420 40.980 442.790 50.080 ;
        RECT 443.365 42.045 443.655 53.880 ;
        RECT 446.815 52.320 447.225 55.415 ;
        RECT 451.270 51.775 451.580 54.290 ;
        RECT 444.260 44.540 444.590 50.735 ;
        RECT 447.180 44.010 447.620 47.285 ;
        RECT 449.560 46.025 450.085 49.965 ;
        RECT 448.720 41.920 449.045 44.685 ;
        RECT 451.235 44.015 451.650 46.405 ;
        RECT 452.265 42.575 452.580 53.260 ;
        RECT 453.595 46.965 454.080 49.975 ;
        RECT 454.775 42.590 455.105 53.285 ;
        RECT 452.965 41.185 453.300 42.535 ;
        RECT 364.635 22.360 364.950 33.410 ;
        RECT 368.470 32.705 368.870 35.755 ;
        RECT 373.390 32.615 373.800 35.710 ;
        RECT 377.970 32.590 378.380 35.685 ;
        RECT 366.305 20.510 366.650 22.970 ;
        RECT 383.420 22.845 383.735 33.530 ;
        RECT 388.655 25.560 389.105 29.720 ;
        RECT 390.355 28.540 390.880 28.980 ;
        RECT 273.040 3.840 273.340 10.770 ;
        RECT 273.695 5.200 273.995 9.260 ;
        RECT 274.350 4.440 274.650 10.790 ;
        RECT 275.665 4.470 275.960 11.295 ;
        RECT 279.505 3.840 279.805 10.780 ;
        RECT 280.185 5.185 280.465 9.275 ;
        RECT 281.715 4.415 282.020 10.775 ;
        RECT 282.565 4.415 282.865 11.235 ;
        RECT 284.295 8.215 284.675 8.235 ;
        RECT 284.295 7.855 284.710 8.215 ;
        RECT 284.330 7.835 284.710 7.855 ;
        RECT 284.305 5.810 284.685 6.190 ;
        RECT 389.455 5.400 389.970 27.635 ;
        RECT 391.140 7.615 391.725 28.315 ;
        RECT 392.735 25.185 393.090 39.125 ;
        RECT 456.080 38.495 456.530 48.760 ;
        RECT 394.360 25.975 394.720 37.525 ;
        RECT 457.245 36.955 457.730 45.840 ;
        RECT 464.185 36.230 464.590 48.275 ;
        RECT 466.260 38.130 466.650 49.555 ;
        RECT 469.420 41.970 469.775 53.055 ;
        RECT 473.165 51.695 473.455 53.755 ;
        RECT 475.935 52.295 476.435 55.345 ;
        RECT 480.905 52.205 481.315 55.300 ;
        RECT 479.945 50.545 480.255 50.575 ;
        RECT 470.745 46.825 471.215 49.815 ;
        RECT 473.095 43.840 473.410 46.210 ;
        RECT 474.715 45.885 475.135 49.850 ;
        RECT 471.380 41.130 471.760 42.505 ;
        RECT 473.820 40.100 474.165 42.560 ;
        RECT 475.455 41.780 475.780 44.545 ;
        RECT 476.440 43.815 476.845 47.145 ;
        RECT 479.945 44.445 480.260 50.545 ;
        RECT 481.090 40.840 481.460 49.940 ;
        RECT 482.035 41.905 482.325 53.740 ;
        RECT 485.485 52.180 485.895 55.275 ;
        RECT 489.940 51.635 490.250 54.150 ;
        RECT 494.190 53.335 494.570 53.715 ;
        RECT 496.320 53.335 496.700 53.715 ;
        RECT 482.930 44.400 483.260 50.595 ;
        RECT 485.835 43.870 486.290 47.145 ;
        RECT 488.195 45.885 488.740 49.825 ;
        RECT 492.250 46.825 492.685 49.835 ;
        RECT 487.390 41.780 487.715 44.545 ;
        RECT 489.905 43.875 490.320 46.265 ;
        RECT 493.445 42.450 493.775 53.145 ;
        RECT 494.880 46.785 495.265 52.570 ;
        RECT 491.635 41.045 491.970 42.395 ;
        RECT 495.240 42.030 495.665 46.305 ;
        RECT 496.940 43.795 497.240 50.835 ;
        RECT 498.060 43.190 498.360 50.120 ;
        RECT 499.370 43.790 499.670 50.140 ;
        RECT 493.900 41.120 494.280 41.500 ;
        RECT 496.095 41.105 496.475 41.485 ;
        RECT 499.965 41.045 500.255 50.825 ;
        RECT 500.685 43.820 500.980 50.645 ;
        RECT 501.815 43.280 502.115 50.090 ;
        RECT 502.605 43.875 502.915 53.915 ;
        RECT 511.795 52.160 512.175 52.540 ;
        RECT 503.400 43.805 503.700 50.635 ;
        RECT 504.525 43.190 504.825 50.130 ;
        RECT 505.975 43.065 506.255 46.100 ;
        RECT 506.735 43.765 507.015 50.125 ;
        RECT 507.585 43.765 507.885 50.585 ;
        RECT 508.725 43.020 509.025 50.175 ;
        RECT 509.370 47.210 509.750 47.590 ;
        RECT 509.370 45.155 509.750 45.535 ;
        RECT 511.220 45.035 511.535 49.360 ;
        RECT 511.830 47.110 512.110 48.640 ;
        RECT 512.400 43.795 512.700 50.835 ;
        RECT 513.520 43.190 513.820 50.120 ;
        RECT 514.175 44.550 514.475 48.610 ;
        RECT 514.830 43.790 515.130 50.140 ;
        RECT 511.695 41.985 512.075 42.365 ;
        RECT 515.425 41.580 515.715 50.825 ;
        RECT 516.145 43.820 516.440 50.645 ;
        RECT 517.275 43.280 517.575 50.090 ;
        RECT 518.065 43.875 518.375 52.610 ;
        RECT 518.860 43.805 519.160 50.635 ;
        RECT 519.985 43.190 520.285 50.130 ;
        RECT 520.665 44.535 520.945 48.625 ;
        RECT 521.435 43.065 521.715 46.100 ;
        RECT 522.195 43.765 522.475 50.125 ;
        RECT 523.045 43.765 523.345 50.585 ;
        RECT 524.185 43.020 524.485 50.175 ;
        RECT 526.525 48.790 526.900 56.990 ;
        RECT 528.270 47.985 528.570 58.980 ;
        RECT 529.200 47.100 529.580 57.355 ;
        RECT 530.070 44.945 530.505 58.520 ;
        RECT 585.780 57.680 586.295 67.980 ;
        RECT 587.465 56.575 588.050 67.355 ;
        RECT 589.015 64.825 589.370 78.745 ;
        RECT 652.360 78.115 652.810 88.380 ;
        RECT 590.640 65.730 591.000 77.145 ;
        RECT 653.525 76.575 654.010 85.460 ;
        RECT 660.190 76.310 660.595 87.840 ;
        RECT 662.265 78.210 662.655 89.310 ;
        RECT 665.690 81.690 666.045 92.775 ;
        RECT 669.435 91.415 669.725 93.475 ;
        RECT 672.205 92.015 672.705 95.065 ;
        RECT 677.175 91.925 677.585 95.020 ;
        RECT 676.215 90.265 676.525 90.295 ;
        RECT 667.015 86.545 667.485 89.535 ;
        RECT 669.365 83.560 669.680 85.930 ;
        RECT 670.985 85.605 671.405 89.570 ;
        RECT 667.650 80.850 668.030 82.225 ;
        RECT 670.090 79.820 670.435 82.280 ;
        RECT 671.725 81.500 672.050 84.265 ;
        RECT 672.710 83.535 673.115 86.865 ;
        RECT 676.215 84.165 676.530 90.265 ;
        RECT 677.360 80.560 677.730 89.660 ;
        RECT 678.305 81.625 678.595 93.460 ;
        RECT 681.755 91.900 682.165 94.995 ;
        RECT 686.210 91.355 686.520 93.870 ;
        RECT 690.460 93.055 690.840 93.435 ;
        RECT 692.590 93.055 692.970 93.435 ;
        RECT 679.200 84.120 679.530 90.315 ;
        RECT 682.105 83.590 682.560 86.865 ;
        RECT 684.465 85.605 685.010 89.545 ;
        RECT 688.520 86.545 688.955 89.555 ;
        RECT 683.660 81.500 683.985 84.265 ;
        RECT 686.175 83.595 686.590 85.985 ;
        RECT 689.715 82.170 690.045 92.865 ;
        RECT 691.150 86.505 691.535 92.290 ;
        RECT 687.905 80.765 688.240 82.115 ;
        RECT 691.510 81.750 691.935 86.025 ;
        RECT 693.210 83.515 693.510 90.555 ;
        RECT 694.330 82.910 694.630 89.840 ;
        RECT 695.640 83.510 695.940 89.860 ;
        RECT 690.170 80.840 690.550 81.220 ;
        RECT 692.365 80.825 692.745 81.205 ;
        RECT 696.235 80.765 696.525 90.545 ;
        RECT 696.955 83.540 697.250 90.365 ;
        RECT 698.085 83.000 698.385 89.810 ;
        RECT 698.875 83.595 699.185 93.635 ;
        RECT 708.065 91.880 708.445 92.260 ;
        RECT 699.670 83.525 699.970 90.355 ;
        RECT 700.795 82.910 701.095 89.850 ;
        RECT 702.245 82.785 702.525 85.820 ;
        RECT 703.005 83.485 703.285 89.845 ;
        RECT 703.855 83.485 704.155 90.305 ;
        RECT 704.995 82.740 705.295 89.895 ;
        RECT 705.640 86.930 706.020 87.310 ;
        RECT 705.640 84.875 706.020 85.255 ;
        RECT 707.490 84.755 707.805 89.080 ;
        RECT 708.100 86.830 708.380 88.360 ;
        RECT 708.670 83.515 708.970 90.555 ;
        RECT 709.790 82.910 710.090 89.840 ;
        RECT 710.445 84.270 710.745 88.330 ;
        RECT 711.100 83.510 711.400 89.860 ;
        RECT 707.965 81.705 708.345 82.085 ;
        RECT 711.695 81.300 711.985 90.545 ;
        RECT 712.415 83.540 712.710 90.365 ;
        RECT 713.545 83.000 713.845 89.810 ;
        RECT 714.335 83.595 714.645 92.330 ;
        RECT 715.130 83.525 715.430 90.355 ;
        RECT 716.255 82.910 716.555 89.850 ;
        RECT 716.935 84.255 717.215 88.345 ;
        RECT 717.705 82.785 717.985 85.820 ;
        RECT 718.465 83.485 718.745 89.845 ;
        RECT 719.315 83.485 719.615 90.305 ;
        RECT 720.455 82.740 720.755 89.895 ;
        RECT 722.740 88.600 723.115 96.885 ;
        RECT 724.485 87.880 724.785 98.875 ;
        RECT 725.565 86.790 725.945 97.045 ;
        RECT 726.435 84.635 726.870 98.210 ;
        RECT 782.140 97.410 782.655 107.460 ;
        RECT 783.825 96.055 784.410 106.835 ;
        RECT 785.705 104.375 786.060 118.165 ;
        RECT 849.050 117.535 849.500 128.035 ;
        RECT 787.330 105.230 787.690 116.565 ;
        RECT 850.215 115.995 850.700 125.235 ;
        RECT 856.630 115.750 857.035 127.280 ;
        RECT 858.705 117.650 859.095 128.750 ;
        RECT 862.110 121.240 862.465 132.325 ;
        RECT 865.855 130.965 866.145 133.025 ;
        RECT 868.625 131.565 869.125 134.615 ;
        RECT 873.595 131.475 874.005 134.570 ;
        RECT 872.635 129.815 872.945 129.845 ;
        RECT 863.435 126.095 863.905 129.085 ;
        RECT 865.785 123.110 866.100 125.480 ;
        RECT 867.405 125.155 867.825 129.120 ;
        RECT 864.070 120.400 864.450 121.775 ;
        RECT 866.510 119.370 866.855 121.830 ;
        RECT 868.145 121.050 868.470 123.815 ;
        RECT 869.130 123.085 869.535 126.415 ;
        RECT 872.635 123.715 872.950 129.815 ;
        RECT 873.780 120.110 874.150 129.210 ;
        RECT 874.725 121.175 875.015 133.010 ;
        RECT 878.175 131.450 878.585 134.545 ;
        RECT 882.630 130.905 882.940 133.420 ;
        RECT 886.880 132.605 887.260 132.985 ;
        RECT 889.010 132.605 889.390 132.985 ;
        RECT 875.620 123.670 875.950 129.865 ;
        RECT 878.525 123.140 878.980 126.415 ;
        RECT 880.885 125.155 881.430 129.095 ;
        RECT 884.940 126.095 885.375 129.105 ;
        RECT 880.080 121.050 880.405 123.815 ;
        RECT 882.595 123.145 883.010 125.535 ;
        RECT 886.135 121.720 886.465 132.415 ;
        RECT 887.570 126.055 887.955 131.840 ;
        RECT 884.325 120.315 884.660 121.665 ;
        RECT 887.930 121.300 888.355 125.575 ;
        RECT 889.630 123.065 889.930 130.105 ;
        RECT 890.750 122.460 891.050 129.390 ;
        RECT 892.060 123.060 892.360 129.410 ;
        RECT 886.590 120.390 886.970 120.770 ;
        RECT 888.785 120.375 889.165 120.755 ;
        RECT 892.655 120.315 892.945 130.095 ;
        RECT 893.375 123.090 893.670 129.915 ;
        RECT 894.505 122.550 894.805 129.360 ;
        RECT 895.295 123.145 895.605 133.185 ;
        RECT 904.485 131.430 904.865 131.810 ;
        RECT 896.090 123.075 896.390 129.905 ;
        RECT 897.215 122.460 897.515 129.400 ;
        RECT 898.665 122.335 898.945 125.370 ;
        RECT 899.425 123.035 899.705 129.395 ;
        RECT 900.275 123.035 900.575 129.855 ;
        RECT 901.415 122.290 901.715 129.445 ;
        RECT 902.060 126.480 902.440 126.860 ;
        RECT 902.060 124.425 902.440 124.805 ;
        RECT 903.910 124.305 904.225 128.630 ;
        RECT 904.520 126.380 904.800 127.910 ;
        RECT 905.090 123.065 905.390 130.105 ;
        RECT 906.210 122.460 906.510 129.390 ;
        RECT 906.865 123.820 907.165 127.880 ;
        RECT 907.520 123.060 907.820 129.410 ;
        RECT 904.385 121.255 904.765 121.635 ;
        RECT 908.115 120.850 908.405 130.095 ;
        RECT 908.835 123.090 909.130 129.915 ;
        RECT 909.965 122.550 910.265 129.360 ;
        RECT 910.755 123.145 911.065 131.880 ;
        RECT 911.550 123.075 911.850 129.905 ;
        RECT 912.675 122.460 912.975 129.400 ;
        RECT 913.355 123.805 913.635 127.895 ;
        RECT 914.125 122.335 914.405 125.370 ;
        RECT 914.885 123.035 915.165 129.395 ;
        RECT 915.735 123.035 916.035 129.855 ;
        RECT 916.875 122.290 917.175 129.445 ;
        RECT 919.060 128.080 919.435 136.280 ;
        RECT 920.805 127.275 921.105 138.270 ;
        RECT 921.950 126.325 922.330 136.580 ;
        RECT 922.820 124.170 923.255 137.745 ;
        RECT 978.525 136.945 979.040 146.995 ;
        RECT 980.210 135.590 980.795 146.370 ;
        RECT 981.835 143.915 982.190 157.705 ;
        RECT 1045.180 157.075 1045.630 167.340 ;
        RECT 983.460 144.770 983.820 156.105 ;
        RECT 1046.345 155.535 1046.830 164.420 ;
        RECT 1052.650 155.160 1053.055 166.690 ;
        RECT 1054.725 157.060 1055.115 168.160 ;
        RECT 1058.495 160.610 1058.850 171.695 ;
        RECT 1062.240 170.335 1062.530 172.395 ;
        RECT 1065.010 170.935 1065.510 173.985 ;
        RECT 1069.980 170.845 1070.390 173.940 ;
        RECT 1069.020 169.185 1069.330 169.215 ;
        RECT 1059.820 165.465 1060.290 168.455 ;
        RECT 1062.170 162.480 1062.485 164.850 ;
        RECT 1063.790 164.525 1064.210 168.490 ;
        RECT 1060.455 159.770 1060.835 161.145 ;
        RECT 1062.895 158.740 1063.240 161.200 ;
        RECT 1064.530 160.420 1064.855 163.185 ;
        RECT 1065.515 162.455 1065.920 165.785 ;
        RECT 1069.020 163.085 1069.335 169.185 ;
        RECT 1070.165 159.480 1070.535 168.580 ;
        RECT 1071.110 160.545 1071.400 172.380 ;
        RECT 1074.560 170.820 1074.970 173.915 ;
        RECT 1079.015 170.275 1079.325 172.790 ;
        RECT 1083.265 171.975 1083.645 172.355 ;
        RECT 1085.395 171.975 1085.775 172.355 ;
        RECT 1072.005 163.040 1072.335 169.235 ;
        RECT 1074.910 162.510 1075.365 165.785 ;
        RECT 1077.270 164.525 1077.815 168.465 ;
        RECT 1081.325 165.465 1081.760 168.475 ;
        RECT 1076.465 160.420 1076.790 163.185 ;
        RECT 1078.980 162.515 1079.395 164.905 ;
        RECT 1082.520 161.090 1082.850 171.785 ;
        RECT 1083.955 165.425 1084.340 171.210 ;
        RECT 1080.710 159.685 1081.045 161.035 ;
        RECT 1084.315 160.670 1084.740 164.945 ;
        RECT 1086.015 162.435 1086.315 169.475 ;
        RECT 1087.135 161.830 1087.435 168.760 ;
        RECT 1088.445 162.430 1088.745 168.780 ;
        RECT 1082.975 159.760 1083.355 160.140 ;
        RECT 1085.170 159.745 1085.550 160.125 ;
        RECT 1089.040 159.685 1089.330 169.465 ;
        RECT 1089.760 162.460 1090.055 169.285 ;
        RECT 1090.890 161.920 1091.190 168.730 ;
        RECT 1091.680 162.515 1091.990 172.555 ;
        RECT 1100.870 170.800 1101.250 171.180 ;
        RECT 1092.475 162.445 1092.775 169.275 ;
        RECT 1093.600 161.830 1093.900 168.770 ;
        RECT 1095.050 161.705 1095.330 164.740 ;
        RECT 1095.810 162.405 1096.090 168.765 ;
        RECT 1096.660 162.405 1096.960 169.225 ;
        RECT 1097.800 161.660 1098.100 168.815 ;
        RECT 1098.445 165.850 1098.825 166.230 ;
        RECT 1098.445 163.795 1098.825 164.175 ;
        RECT 1100.295 163.675 1100.610 168.000 ;
        RECT 1100.905 165.750 1101.185 167.280 ;
        RECT 1101.475 162.435 1101.775 169.475 ;
        RECT 1103.250 163.190 1103.550 167.250 ;
        RECT 1100.770 160.625 1101.150 161.005 ;
        RECT 1104.500 160.220 1104.790 169.465 ;
        RECT 1106.350 161.920 1106.650 168.730 ;
        RECT 1107.140 162.515 1107.450 171.250 ;
        RECT 1107.935 162.445 1108.235 169.275 ;
        RECT 1109.740 163.175 1110.020 167.265 ;
        RECT 1110.510 161.705 1110.790 164.740 ;
        RECT 1113.260 161.660 1113.560 168.815 ;
        RECT 1150.120 160.695 1150.435 171.745 ;
        RECT 1153.955 171.040 1154.355 174.090 ;
        RECT 1158.875 170.950 1159.285 174.045 ;
        RECT 1163.455 170.925 1163.865 174.020 ;
        RECT 1151.790 158.845 1152.135 161.305 ;
        RECT 1168.905 161.180 1169.220 171.865 ;
        RECT 1174.090 163.970 1174.540 168.130 ;
        RECT 1183.495 167.670 1183.875 168.050 ;
        RECT 1175.790 166.950 1176.315 167.390 ;
        RECT 1183.485 166.920 1183.865 167.300 ;
        RECT 987.110 147.980 987.490 148.360 ;
        RECT 987.100 147.230 987.480 147.610 ;
        RECT 987.145 146.545 987.525 146.925 ;
        RECT 987.110 145.875 987.490 146.255 ;
        RECT 987.825 142.800 988.125 149.840 ;
        RECT 988.945 142.195 989.245 149.125 ;
        RECT 989.600 143.555 989.900 147.615 ;
        RECT 990.255 142.795 990.555 149.145 ;
        RECT 990.850 144.670 991.170 149.830 ;
        RECT 991.570 142.825 991.865 149.650 ;
        RECT 992.700 142.285 993.000 149.095 ;
        RECT 993.490 142.880 993.800 149.070 ;
        RECT 994.285 142.810 994.585 149.640 ;
        RECT 995.410 142.195 995.710 149.135 ;
        RECT 996.090 143.540 996.370 147.630 ;
        RECT 996.860 142.070 997.140 145.105 ;
        RECT 997.620 142.770 997.925 149.130 ;
        RECT 998.470 142.770 998.770 149.590 ;
        RECT 999.610 142.025 999.910 149.180 ;
        RECT 1000.275 147.980 1000.655 148.360 ;
        RECT 1002.545 147.980 1002.925 148.385 ;
        RECT 1000.280 147.230 1000.660 147.610 ;
        RECT 1002.550 147.230 1002.930 147.635 ;
        RECT 1000.280 146.215 1000.660 146.595 ;
        RECT 1002.065 144.795 1002.385 146.925 ;
        RECT 1000.495 141.505 1000.875 144.525 ;
        RECT 1002.675 143.955 1002.955 146.360 ;
        RECT 1003.285 142.800 1003.585 149.840 ;
        RECT 1004.405 142.195 1004.705 149.125 ;
        RECT 1005.060 143.555 1005.360 147.615 ;
        RECT 1005.715 142.795 1006.015 149.145 ;
        RECT 1006.310 144.670 1006.635 149.830 ;
        RECT 1007.030 142.825 1007.325 149.650 ;
        RECT 1008.160 142.285 1008.460 149.095 ;
        RECT 1008.950 142.880 1009.260 149.070 ;
        RECT 1009.745 142.810 1010.045 149.640 ;
        RECT 1010.870 142.195 1011.170 149.135 ;
        RECT 1011.550 143.540 1011.830 147.630 ;
        RECT 1012.320 142.070 1012.600 145.105 ;
        RECT 1013.080 142.770 1013.400 149.130 ;
        RECT 1013.930 142.770 1014.230 149.590 ;
        RECT 1015.070 142.025 1015.370 149.180 ;
        RECT 1016.010 147.980 1016.370 149.810 ;
        RECT 1015.705 144.170 1016.085 144.550 ;
        RECT 1016.410 140.055 1016.770 146.615 ;
        RECT 1017.550 144.805 1017.875 146.670 ;
        RECT 1018.190 146.460 1018.605 149.810 ;
        RECT 1018.215 141.460 1018.675 146.145 ;
        RECT 1019.000 144.005 1019.450 152.825 ;
        RECT 1019.860 141.630 1020.215 151.935 ;
        RECT 1020.525 147.235 1020.870 148.290 ;
        RECT 1021.185 145.830 1021.615 148.820 ;
        RECT 1018.930 140.115 1019.310 140.495 ;
        RECT 1021.820 140.135 1022.200 141.510 ;
        RECT 1022.590 140.955 1022.905 152.005 ;
        RECT 1023.605 150.700 1023.895 152.760 ;
        RECT 1026.390 151.300 1026.865 154.350 ;
        RECT 1031.345 151.210 1031.755 154.305 ;
        RECT 1030.385 149.550 1030.695 149.580 ;
        RECT 1023.525 142.845 1023.850 145.215 ;
        RECT 1025.175 144.890 1025.575 148.855 ;
        RECT 1024.260 139.105 1024.605 141.565 ;
        RECT 1025.895 140.785 1026.220 143.550 ;
        RECT 1026.880 142.820 1027.285 146.150 ;
        RECT 1030.385 143.450 1030.700 149.550 ;
        RECT 1031.530 139.845 1031.900 148.945 ;
        RECT 1032.475 140.910 1032.765 152.745 ;
        RECT 1035.925 151.185 1036.335 154.280 ;
        RECT 1040.380 150.640 1040.690 153.155 ;
        RECT 1033.370 143.405 1033.700 149.600 ;
        RECT 1036.290 142.875 1036.730 146.150 ;
        RECT 1038.670 144.890 1039.195 148.830 ;
        RECT 1037.830 140.785 1038.155 143.550 ;
        RECT 1040.345 142.880 1040.760 145.270 ;
        RECT 1041.375 141.440 1041.690 152.125 ;
        RECT 1042.705 145.830 1043.190 148.840 ;
        RECT 1043.885 141.455 1044.215 152.150 ;
        RECT 1042.075 140.050 1042.410 141.400 ;
        RECT 953.770 121.170 954.085 132.220 ;
        RECT 957.605 131.515 958.005 134.565 ;
        RECT 962.525 131.425 962.935 134.520 ;
        RECT 967.105 131.400 967.515 134.495 ;
        RECT 955.440 119.320 955.785 121.780 ;
        RECT 972.555 121.655 972.870 132.340 ;
        RECT 977.740 124.445 978.190 128.605 ;
        RECT 979.440 127.425 979.965 127.865 ;
        RECT 790.765 108.430 791.145 108.810 ;
        RECT 790.755 107.680 791.135 108.060 ;
        RECT 790.800 106.995 791.180 107.375 ;
        RECT 790.765 106.325 791.145 106.705 ;
        RECT 791.480 103.250 791.780 110.290 ;
        RECT 792.600 102.645 792.900 109.575 ;
        RECT 793.255 104.005 793.555 108.065 ;
        RECT 793.910 103.245 794.210 109.595 ;
        RECT 794.505 105.120 794.825 110.280 ;
        RECT 795.225 103.275 795.520 110.100 ;
        RECT 796.355 102.735 796.655 109.545 ;
        RECT 797.145 103.330 797.455 109.520 ;
        RECT 797.940 103.260 798.240 110.090 ;
        RECT 799.065 102.645 799.365 109.585 ;
        RECT 799.745 103.990 800.025 108.080 ;
        RECT 800.515 102.520 800.795 105.555 ;
        RECT 801.275 103.220 801.580 109.580 ;
        RECT 802.125 103.220 802.425 110.040 ;
        RECT 803.265 102.475 803.565 109.630 ;
        RECT 803.930 108.430 804.310 108.810 ;
        RECT 806.200 108.430 806.580 108.835 ;
        RECT 803.935 107.680 804.315 108.060 ;
        RECT 806.205 107.680 806.585 108.085 ;
        RECT 803.935 106.665 804.315 107.045 ;
        RECT 805.720 105.245 806.040 107.375 ;
        RECT 804.150 101.955 804.530 104.975 ;
        RECT 806.330 104.405 806.610 106.810 ;
        RECT 806.940 103.250 807.240 110.290 ;
        RECT 808.060 102.645 808.360 109.575 ;
        RECT 808.715 104.005 809.015 108.065 ;
        RECT 809.370 103.245 809.670 109.595 ;
        RECT 809.965 105.120 810.290 110.280 ;
        RECT 810.685 103.275 810.980 110.100 ;
        RECT 811.815 102.735 812.115 109.545 ;
        RECT 812.605 103.330 812.915 109.520 ;
        RECT 813.400 103.260 813.700 110.090 ;
        RECT 814.525 102.645 814.825 109.585 ;
        RECT 815.205 103.990 815.485 108.080 ;
        RECT 815.975 102.520 816.255 105.555 ;
        RECT 816.735 103.220 817.055 109.580 ;
        RECT 817.585 103.220 817.885 110.040 ;
        RECT 818.725 102.475 819.025 109.630 ;
        RECT 819.665 108.430 820.025 110.260 ;
        RECT 819.360 104.620 819.740 105.000 ;
        RECT 820.065 100.505 820.425 107.065 ;
        RECT 821.205 105.255 821.530 107.120 ;
        RECT 821.845 106.910 822.260 110.260 ;
        RECT 821.870 101.910 822.330 106.595 ;
        RECT 822.655 104.455 823.105 113.275 ;
        RECT 823.515 102.080 823.870 112.385 ;
        RECT 824.180 107.685 824.525 108.740 ;
        RECT 824.840 106.280 825.270 109.270 ;
        RECT 822.585 100.565 822.965 100.945 ;
        RECT 825.475 100.585 825.855 101.960 ;
        RECT 826.245 101.405 826.560 112.455 ;
        RECT 827.260 111.150 827.550 113.210 ;
        RECT 830.045 111.750 830.520 114.800 ;
        RECT 835.000 111.660 835.410 114.755 ;
        RECT 834.040 110.000 834.350 110.030 ;
        RECT 827.180 103.295 827.505 105.665 ;
        RECT 828.830 105.340 829.230 109.305 ;
        RECT 827.915 99.555 828.260 102.015 ;
        RECT 829.550 101.235 829.875 104.000 ;
        RECT 830.535 103.270 830.940 106.600 ;
        RECT 834.040 103.900 834.355 110.000 ;
        RECT 835.185 100.295 835.555 109.395 ;
        RECT 836.130 101.360 836.420 113.195 ;
        RECT 839.580 111.635 839.990 114.730 ;
        RECT 844.035 111.090 844.345 113.605 ;
        RECT 837.025 103.855 837.355 110.050 ;
        RECT 839.945 103.325 840.385 106.600 ;
        RECT 842.325 105.340 842.850 109.280 ;
        RECT 841.485 101.235 841.810 104.000 ;
        RECT 844.000 103.330 844.415 105.720 ;
        RECT 845.030 101.890 845.345 112.575 ;
        RECT 846.360 106.280 846.845 109.290 ;
        RECT 847.540 101.905 847.870 112.600 ;
        RECT 845.730 100.500 846.065 101.850 ;
        RECT 757.345 81.690 757.660 92.740 ;
        RECT 761.180 92.035 761.580 95.085 ;
        RECT 766.100 91.945 766.510 95.040 ;
        RECT 770.680 91.920 771.090 95.015 ;
        RECT 759.015 79.840 759.360 82.300 ;
        RECT 776.130 82.175 776.445 92.860 ;
        RECT 781.315 84.965 781.765 89.125 ;
        RECT 783.015 87.945 783.540 88.385 ;
        RECT 594.425 68.960 594.805 69.340 ;
        RECT 594.415 68.210 594.795 68.590 ;
        RECT 594.460 67.525 594.840 67.905 ;
        RECT 594.425 66.855 594.805 67.235 ;
        RECT 595.140 63.780 595.440 70.820 ;
        RECT 596.260 63.175 596.560 70.105 ;
        RECT 596.915 64.535 597.215 68.595 ;
        RECT 597.570 63.775 597.870 70.125 ;
        RECT 598.165 65.650 598.485 70.810 ;
        RECT 598.885 63.805 599.180 70.630 ;
        RECT 600.015 63.265 600.315 70.075 ;
        RECT 600.805 63.860 601.115 70.050 ;
        RECT 601.600 63.790 601.900 70.620 ;
        RECT 602.725 63.175 603.025 70.115 ;
        RECT 603.405 64.520 603.685 68.610 ;
        RECT 604.175 63.050 604.455 66.085 ;
        RECT 604.935 63.750 605.240 70.110 ;
        RECT 605.785 63.750 606.085 70.570 ;
        RECT 606.925 63.005 607.225 70.160 ;
        RECT 607.590 68.960 607.970 69.340 ;
        RECT 609.860 68.960 610.240 69.365 ;
        RECT 607.595 68.210 607.975 68.590 ;
        RECT 609.865 68.210 610.245 68.615 ;
        RECT 607.595 67.195 607.975 67.575 ;
        RECT 609.380 65.775 609.700 67.905 ;
        RECT 607.810 62.485 608.190 65.505 ;
        RECT 609.990 64.935 610.270 67.340 ;
        RECT 610.600 63.780 610.900 70.820 ;
        RECT 611.720 63.175 612.020 70.105 ;
        RECT 612.375 64.535 612.675 68.595 ;
        RECT 613.030 63.775 613.330 70.125 ;
        RECT 613.625 65.650 613.950 70.810 ;
        RECT 614.345 63.805 614.640 70.630 ;
        RECT 615.475 63.265 615.775 70.075 ;
        RECT 616.265 63.860 616.575 70.050 ;
        RECT 617.060 63.790 617.360 70.620 ;
        RECT 618.185 63.175 618.485 70.115 ;
        RECT 618.865 64.520 619.145 68.610 ;
        RECT 619.635 63.050 619.915 66.085 ;
        RECT 620.395 63.750 620.715 70.110 ;
        RECT 621.245 63.750 621.545 70.570 ;
        RECT 622.385 63.005 622.685 70.160 ;
        RECT 623.325 68.960 623.685 70.790 ;
        RECT 623.020 65.150 623.400 65.530 ;
        RECT 623.725 61.035 624.085 67.595 ;
        RECT 624.865 65.785 625.190 67.650 ;
        RECT 625.505 67.440 625.920 70.790 ;
        RECT 625.530 62.440 625.990 67.125 ;
        RECT 626.315 64.985 626.765 73.805 ;
        RECT 627.175 62.610 627.530 72.915 ;
        RECT 627.840 68.215 628.185 69.270 ;
        RECT 628.500 66.810 628.930 69.800 ;
        RECT 626.245 61.095 626.625 61.475 ;
        RECT 629.135 61.115 629.515 62.490 ;
        RECT 629.905 61.935 630.220 72.985 ;
        RECT 630.920 71.680 631.210 73.740 ;
        RECT 633.705 72.280 634.180 75.330 ;
        RECT 638.660 72.190 639.070 75.285 ;
        RECT 637.700 70.530 638.010 70.560 ;
        RECT 630.840 63.825 631.165 66.195 ;
        RECT 632.490 65.870 632.890 69.835 ;
        RECT 631.575 60.085 631.920 62.545 ;
        RECT 633.210 61.765 633.535 64.530 ;
        RECT 634.195 63.800 634.600 67.130 ;
        RECT 637.700 64.430 638.015 70.530 ;
        RECT 638.845 60.825 639.215 69.925 ;
        RECT 639.790 61.890 640.080 73.725 ;
        RECT 643.240 72.165 643.650 75.260 ;
        RECT 647.695 71.620 648.005 74.135 ;
        RECT 640.685 64.385 641.015 70.580 ;
        RECT 643.605 63.855 644.045 67.130 ;
        RECT 645.985 65.870 646.510 69.810 ;
        RECT 645.145 61.765 645.470 64.530 ;
        RECT 647.660 63.860 648.075 66.250 ;
        RECT 648.690 62.420 649.005 73.105 ;
        RECT 650.020 66.810 650.505 69.820 ;
        RECT 651.200 62.435 651.530 73.130 ;
        RECT 649.390 61.030 649.725 62.380 ;
        RECT 560.980 42.135 561.295 53.185 ;
        RECT 564.815 52.480 565.215 55.530 ;
        RECT 569.735 52.390 570.145 55.485 ;
        RECT 574.315 52.365 574.725 55.460 ;
        RECT 562.650 40.285 562.995 42.745 ;
        RECT 579.765 42.620 580.080 53.305 ;
        RECT 584.950 45.410 585.400 49.570 ;
        RECT 586.650 48.390 587.175 48.830 ;
        RECT 397.970 29.320 398.350 29.700 ;
        RECT 397.960 28.570 398.340 28.950 ;
        RECT 398.005 27.885 398.385 28.265 ;
        RECT 397.970 27.215 398.350 27.595 ;
        RECT 398.685 24.140 398.985 31.180 ;
        RECT 399.805 23.535 400.105 30.465 ;
        RECT 400.460 24.895 400.760 28.955 ;
        RECT 401.115 24.135 401.415 30.485 ;
        RECT 401.710 26.010 402.030 31.170 ;
        RECT 402.430 24.165 402.725 30.990 ;
        RECT 403.560 23.625 403.860 30.435 ;
        RECT 404.350 24.220 404.660 30.410 ;
        RECT 405.145 24.150 405.445 30.980 ;
        RECT 406.270 23.535 406.570 30.475 ;
        RECT 406.950 24.880 407.230 28.970 ;
        RECT 407.720 23.410 408.000 26.445 ;
        RECT 408.480 24.110 408.785 30.470 ;
        RECT 409.330 24.110 409.630 30.930 ;
        RECT 410.470 23.365 410.770 30.520 ;
        RECT 411.135 29.320 411.515 29.700 ;
        RECT 413.405 29.320 413.785 29.725 ;
        RECT 411.140 28.570 411.520 28.950 ;
        RECT 413.410 28.570 413.790 28.975 ;
        RECT 411.140 27.555 411.520 27.935 ;
        RECT 412.925 26.135 413.245 28.265 ;
        RECT 411.355 22.845 411.735 25.865 ;
        RECT 413.535 25.295 413.815 27.700 ;
        RECT 414.145 24.140 414.445 31.180 ;
        RECT 415.265 23.535 415.565 30.465 ;
        RECT 415.920 24.895 416.220 28.955 ;
        RECT 416.575 24.135 416.875 30.485 ;
        RECT 417.170 26.010 417.495 31.170 ;
        RECT 417.890 24.165 418.185 30.990 ;
        RECT 419.020 23.625 419.320 30.435 ;
        RECT 419.810 24.220 420.120 30.410 ;
        RECT 420.605 24.150 420.905 30.980 ;
        RECT 421.730 23.535 422.030 30.475 ;
        RECT 422.410 24.880 422.690 28.970 ;
        RECT 423.180 23.410 423.460 26.445 ;
        RECT 423.940 24.110 424.260 30.470 ;
        RECT 424.790 24.110 425.090 30.930 ;
        RECT 425.930 23.365 426.230 30.520 ;
        RECT 426.870 29.320 427.230 31.150 ;
        RECT 426.565 25.510 426.945 25.890 ;
        RECT 427.270 21.395 427.630 27.955 ;
        RECT 428.410 26.145 428.735 28.010 ;
        RECT 429.050 27.800 429.465 31.150 ;
        RECT 429.075 22.800 429.535 27.485 ;
        RECT 429.860 25.345 430.310 34.165 ;
        RECT 430.720 22.970 431.075 33.275 ;
        RECT 431.385 28.575 431.730 29.630 ;
        RECT 432.045 27.170 432.475 30.160 ;
        RECT 429.790 21.455 430.170 21.835 ;
        RECT 432.680 21.475 433.060 22.850 ;
        RECT 433.450 22.295 433.765 33.345 ;
        RECT 434.465 32.040 434.755 34.100 ;
        RECT 437.250 32.640 437.725 35.690 ;
        RECT 442.205 32.550 442.615 35.645 ;
        RECT 441.245 30.890 441.555 30.920 ;
        RECT 434.385 24.185 434.710 26.555 ;
        RECT 436.035 26.230 436.435 30.195 ;
        RECT 435.120 20.445 435.465 22.905 ;
        RECT 436.755 22.125 437.080 24.890 ;
        RECT 437.740 24.160 438.145 27.490 ;
        RECT 441.245 24.790 441.560 30.890 ;
        RECT 442.390 21.185 442.760 30.285 ;
        RECT 443.335 22.250 443.625 34.085 ;
        RECT 446.785 32.525 447.195 35.620 ;
        RECT 451.240 31.980 451.550 34.495 ;
        RECT 444.230 24.745 444.560 30.940 ;
        RECT 447.150 24.215 447.590 27.490 ;
        RECT 449.530 26.230 450.055 30.170 ;
        RECT 448.690 22.125 449.015 24.890 ;
        RECT 451.205 24.220 451.620 26.610 ;
        RECT 452.235 22.780 452.550 33.465 ;
        RECT 453.565 27.170 454.050 30.180 ;
        RECT 454.745 22.795 455.075 33.490 ;
        RECT 460.025 29.090 463.350 29.680 ;
        RECT 460.025 28.475 460.775 29.090 ;
        RECT 461.930 25.635 462.600 28.285 ;
        RECT 452.935 21.390 453.270 22.740 ;
        RECT 463.890 9.480 464.340 28.520 ;
        RECT 465.680 8.705 466.095 29.885 ;
        RECT 469.420 22.305 469.775 33.390 ;
        RECT 473.165 32.030 473.455 34.090 ;
        RECT 475.935 32.630 476.435 35.680 ;
        RECT 480.905 32.540 481.315 35.635 ;
        RECT 479.945 30.880 480.255 30.910 ;
        RECT 470.745 27.160 471.215 30.150 ;
        RECT 473.095 24.175 473.410 26.545 ;
        RECT 474.715 26.220 475.135 30.185 ;
        RECT 471.380 21.465 471.760 22.840 ;
        RECT 473.820 20.435 474.165 22.895 ;
        RECT 475.455 22.115 475.780 24.880 ;
        RECT 476.440 24.150 476.845 27.480 ;
        RECT 479.945 24.780 480.260 30.880 ;
        RECT 481.090 21.175 481.460 30.275 ;
        RECT 482.035 22.240 482.325 34.075 ;
        RECT 485.485 32.515 485.895 35.610 ;
        RECT 489.940 31.970 490.250 34.485 ;
        RECT 494.190 33.670 494.570 34.050 ;
        RECT 496.320 33.670 496.700 34.050 ;
        RECT 482.930 24.735 483.260 30.930 ;
        RECT 485.835 24.205 486.290 27.480 ;
        RECT 488.195 26.220 488.740 30.160 ;
        RECT 492.250 27.160 492.685 30.170 ;
        RECT 487.390 22.115 487.715 24.880 ;
        RECT 489.905 24.210 490.320 26.600 ;
        RECT 493.445 22.785 493.775 33.480 ;
        RECT 494.880 27.120 495.265 32.905 ;
        RECT 491.635 21.380 491.970 22.730 ;
        RECT 495.240 22.365 495.665 26.640 ;
        RECT 496.940 24.130 497.240 31.170 ;
        RECT 498.060 23.525 498.360 30.455 ;
        RECT 499.370 24.125 499.670 30.475 ;
        RECT 493.900 21.455 494.280 21.835 ;
        RECT 496.095 21.440 496.475 21.820 ;
        RECT 499.965 21.380 500.255 31.160 ;
        RECT 500.685 24.155 500.980 30.980 ;
        RECT 501.815 23.615 502.115 30.425 ;
        RECT 502.605 24.210 502.915 34.250 ;
        RECT 511.795 32.495 512.175 32.875 ;
        RECT 503.400 24.140 503.700 30.970 ;
        RECT 504.525 23.525 504.825 30.465 ;
        RECT 505.975 23.400 506.255 26.435 ;
        RECT 506.735 24.100 507.015 30.460 ;
        RECT 507.585 24.100 507.885 30.920 ;
        RECT 508.725 23.355 509.025 30.510 ;
        RECT 509.370 27.545 509.750 27.925 ;
        RECT 509.370 25.490 509.750 25.870 ;
        RECT 511.220 25.370 511.535 29.695 ;
        RECT 511.830 27.445 512.110 28.975 ;
        RECT 512.400 24.130 512.700 31.170 ;
        RECT 513.520 23.525 513.820 30.455 ;
        RECT 514.175 24.885 514.475 28.945 ;
        RECT 514.830 24.125 515.130 30.475 ;
        RECT 511.695 22.320 512.075 22.700 ;
        RECT 515.425 21.915 515.715 31.160 ;
        RECT 516.145 24.155 516.440 30.980 ;
        RECT 517.275 23.615 517.575 30.425 ;
        RECT 518.065 24.210 518.375 32.945 ;
        RECT 518.860 24.140 519.160 30.970 ;
        RECT 519.985 23.525 520.285 30.465 ;
        RECT 520.665 24.870 520.945 28.960 ;
        RECT 521.435 23.400 521.715 26.435 ;
        RECT 522.195 24.100 522.475 30.460 ;
        RECT 523.045 24.100 523.345 30.920 ;
        RECT 524.185 23.355 524.485 30.510 ;
        RECT 526.110 29.275 526.485 37.115 ;
        RECT 527.965 28.525 528.265 39.065 ;
        RECT 529.200 27.440 529.580 37.695 ;
        RECT 530.070 25.285 530.505 38.860 ;
        RECT 585.780 38.125 586.295 48.175 ;
        RECT 587.465 36.770 588.050 47.550 ;
        RECT 589.110 45.060 589.465 58.970 ;
        RECT 652.455 58.340 652.905 68.605 ;
        RECT 590.735 45.980 591.095 57.370 ;
        RECT 653.620 56.800 654.105 65.685 ;
        RECT 660.450 56.155 660.855 68.035 ;
        RECT 662.525 58.055 662.915 69.635 ;
        RECT 665.795 61.975 666.150 73.060 ;
        RECT 669.540 71.700 669.830 73.760 ;
        RECT 672.310 72.300 672.810 75.350 ;
        RECT 677.280 72.210 677.690 75.305 ;
        RECT 676.320 70.550 676.630 70.580 ;
        RECT 667.120 66.830 667.590 69.820 ;
        RECT 669.470 63.845 669.785 66.215 ;
        RECT 671.090 65.890 671.510 69.855 ;
        RECT 667.755 61.135 668.135 62.510 ;
        RECT 670.195 60.105 670.540 62.565 ;
        RECT 671.830 61.785 672.155 64.550 ;
        RECT 672.815 63.820 673.220 67.150 ;
        RECT 676.320 64.450 676.635 70.550 ;
        RECT 677.465 60.845 677.835 69.945 ;
        RECT 678.410 61.910 678.700 73.745 ;
        RECT 681.860 72.185 682.270 75.280 ;
        RECT 686.315 71.640 686.625 74.155 ;
        RECT 690.565 73.340 690.945 73.720 ;
        RECT 692.695 73.340 693.075 73.720 ;
        RECT 679.305 64.405 679.635 70.600 ;
        RECT 682.210 63.875 682.665 67.150 ;
        RECT 684.570 65.890 685.115 69.830 ;
        RECT 688.625 66.830 689.060 69.840 ;
        RECT 683.765 61.785 684.090 64.550 ;
        RECT 686.280 63.880 686.695 66.270 ;
        RECT 689.820 62.455 690.150 73.150 ;
        RECT 691.255 66.790 691.640 72.575 ;
        RECT 688.010 61.050 688.345 62.400 ;
        RECT 691.615 62.035 692.040 66.310 ;
        RECT 693.315 63.800 693.615 70.840 ;
        RECT 694.435 63.195 694.735 70.125 ;
        RECT 695.745 63.795 696.045 70.145 ;
        RECT 690.275 61.125 690.655 61.505 ;
        RECT 692.470 61.110 692.850 61.490 ;
        RECT 696.340 61.050 696.630 70.830 ;
        RECT 697.060 63.825 697.355 70.650 ;
        RECT 698.190 63.285 698.490 70.095 ;
        RECT 698.980 63.880 699.290 73.920 ;
        RECT 708.170 72.165 708.550 72.545 ;
        RECT 699.775 63.810 700.075 70.640 ;
        RECT 700.900 63.195 701.200 70.135 ;
        RECT 702.350 63.070 702.630 66.105 ;
        RECT 703.110 63.770 703.390 70.130 ;
        RECT 703.960 63.770 704.260 70.590 ;
        RECT 705.100 63.025 705.400 70.180 ;
        RECT 705.745 67.215 706.125 67.595 ;
        RECT 705.745 65.160 706.125 65.540 ;
        RECT 707.595 65.040 707.910 69.365 ;
        RECT 708.205 67.115 708.485 68.645 ;
        RECT 708.775 63.800 709.075 70.840 ;
        RECT 709.895 63.195 710.195 70.125 ;
        RECT 710.550 64.555 710.850 68.615 ;
        RECT 711.205 63.795 711.505 70.145 ;
        RECT 708.070 61.990 708.450 62.370 ;
        RECT 711.800 61.585 712.090 70.830 ;
        RECT 712.520 63.825 712.815 70.650 ;
        RECT 713.650 63.285 713.950 70.095 ;
        RECT 714.440 63.880 714.750 72.615 ;
        RECT 715.235 63.810 715.535 70.640 ;
        RECT 716.360 63.195 716.660 70.135 ;
        RECT 717.040 64.540 717.320 68.630 ;
        RECT 717.810 63.070 718.090 66.105 ;
        RECT 718.570 63.770 718.850 70.130 ;
        RECT 719.420 63.770 719.720 70.590 ;
        RECT 720.560 63.025 720.860 70.180 ;
        RECT 722.640 68.900 723.015 77.180 ;
        RECT 724.385 68.060 724.685 79.170 ;
        RECT 725.565 67.080 725.945 77.335 ;
        RECT 726.435 64.925 726.870 78.500 ;
        RECT 782.145 77.700 782.660 87.750 ;
        RECT 783.830 76.345 784.415 87.125 ;
        RECT 785.660 84.585 786.015 98.375 ;
        RECT 849.005 97.745 849.455 108.235 ;
        RECT 787.285 85.490 787.645 96.775 ;
        RECT 850.170 96.205 850.655 105.365 ;
        RECT 856.630 96.015 857.035 107.545 ;
        RECT 858.705 97.915 859.095 109.015 ;
        RECT 862.110 101.445 862.465 112.530 ;
        RECT 865.855 111.170 866.145 113.230 ;
        RECT 868.625 111.770 869.125 114.820 ;
        RECT 873.595 111.680 874.005 114.775 ;
        RECT 872.635 110.020 872.945 110.050 ;
        RECT 863.435 106.300 863.905 109.290 ;
        RECT 865.785 103.315 866.100 105.685 ;
        RECT 867.405 105.360 867.825 109.325 ;
        RECT 864.070 100.605 864.450 101.980 ;
        RECT 866.510 99.575 866.855 102.035 ;
        RECT 868.145 101.255 868.470 104.020 ;
        RECT 869.130 103.290 869.535 106.620 ;
        RECT 872.635 103.920 872.950 110.020 ;
        RECT 873.780 100.315 874.150 109.415 ;
        RECT 874.725 101.380 875.015 113.215 ;
        RECT 878.175 111.655 878.585 114.750 ;
        RECT 882.630 111.110 882.940 113.625 ;
        RECT 886.880 112.810 887.260 113.190 ;
        RECT 889.010 112.810 889.390 113.190 ;
        RECT 875.620 103.875 875.950 110.070 ;
        RECT 878.525 103.345 878.980 106.620 ;
        RECT 880.885 105.360 881.430 109.300 ;
        RECT 884.940 106.300 885.375 109.310 ;
        RECT 880.080 101.255 880.405 104.020 ;
        RECT 882.595 103.350 883.010 105.740 ;
        RECT 886.135 101.925 886.465 112.620 ;
        RECT 887.570 106.260 887.955 112.045 ;
        RECT 884.325 100.520 884.660 101.870 ;
        RECT 887.930 101.505 888.355 105.780 ;
        RECT 889.630 103.270 889.930 110.310 ;
        RECT 890.750 102.665 891.050 109.595 ;
        RECT 892.060 103.265 892.360 109.615 ;
        RECT 886.590 100.595 886.970 100.975 ;
        RECT 888.785 100.580 889.165 100.960 ;
        RECT 892.655 100.520 892.945 110.300 ;
        RECT 893.375 103.295 893.670 110.120 ;
        RECT 894.505 102.755 894.805 109.565 ;
        RECT 895.295 103.350 895.605 113.390 ;
        RECT 904.485 111.635 904.865 112.015 ;
        RECT 896.090 103.280 896.390 110.110 ;
        RECT 897.215 102.665 897.515 109.605 ;
        RECT 898.665 102.540 898.945 105.575 ;
        RECT 899.425 103.240 899.705 109.600 ;
        RECT 900.275 103.240 900.575 110.060 ;
        RECT 901.415 102.495 901.715 109.650 ;
        RECT 902.060 106.685 902.440 107.065 ;
        RECT 902.060 104.630 902.440 105.010 ;
        RECT 903.910 104.510 904.225 108.835 ;
        RECT 904.520 106.585 904.800 108.115 ;
        RECT 905.090 103.270 905.390 110.310 ;
        RECT 906.210 102.665 906.510 109.595 ;
        RECT 906.865 104.025 907.165 108.085 ;
        RECT 907.520 103.265 907.820 109.615 ;
        RECT 904.385 101.460 904.765 101.840 ;
        RECT 908.115 101.055 908.405 110.300 ;
        RECT 908.835 103.295 909.130 110.120 ;
        RECT 909.965 102.755 910.265 109.565 ;
        RECT 910.755 103.350 911.065 112.085 ;
        RECT 911.550 103.280 911.850 110.110 ;
        RECT 912.675 102.665 912.975 109.605 ;
        RECT 913.355 104.010 913.635 108.100 ;
        RECT 914.125 102.540 914.405 105.575 ;
        RECT 914.885 103.240 915.165 109.600 ;
        RECT 915.735 103.240 916.035 110.060 ;
        RECT 916.875 102.495 917.175 109.650 ;
        RECT 919.080 108.420 919.455 116.620 ;
        RECT 920.825 107.615 921.125 118.610 ;
        RECT 921.950 106.530 922.330 116.785 ;
        RECT 922.820 104.375 923.255 117.950 ;
        RECT 978.675 117.230 979.190 127.280 ;
        RECT 980.360 115.875 980.945 126.655 ;
        RECT 981.835 124.150 982.190 138.205 ;
        RECT 1045.180 137.575 1045.630 147.690 ;
        RECT 983.460 124.955 983.820 136.605 ;
        RECT 1046.345 136.035 1046.830 144.790 ;
        RECT 1052.950 135.410 1053.355 146.940 ;
        RECT 1055.025 137.310 1055.415 148.410 ;
        RECT 1058.295 140.885 1058.650 151.970 ;
        RECT 1062.040 150.610 1062.330 152.670 ;
        RECT 1064.810 151.210 1065.310 154.260 ;
        RECT 1069.780 151.120 1070.190 154.215 ;
        RECT 1068.820 149.460 1069.130 149.490 ;
        RECT 1059.620 145.740 1060.090 148.730 ;
        RECT 1061.970 142.755 1062.285 145.125 ;
        RECT 1063.590 144.800 1064.010 148.765 ;
        RECT 1060.255 140.045 1060.635 141.420 ;
        RECT 1062.695 139.015 1063.040 141.475 ;
        RECT 1064.330 140.695 1064.655 143.460 ;
        RECT 1065.315 142.730 1065.720 146.060 ;
        RECT 1068.820 143.360 1069.135 149.460 ;
        RECT 1069.965 139.755 1070.335 148.855 ;
        RECT 1070.910 140.820 1071.200 152.655 ;
        RECT 1074.360 151.095 1074.770 154.190 ;
        RECT 1078.815 150.550 1079.125 153.065 ;
        RECT 1083.065 152.250 1083.445 152.630 ;
        RECT 1085.195 152.250 1085.575 152.630 ;
        RECT 1071.805 143.315 1072.135 149.510 ;
        RECT 1074.710 142.785 1075.165 146.060 ;
        RECT 1077.070 144.800 1077.615 148.740 ;
        RECT 1081.125 145.740 1081.560 148.750 ;
        RECT 1076.265 140.695 1076.590 143.460 ;
        RECT 1078.780 142.790 1079.195 145.180 ;
        RECT 1082.320 141.365 1082.650 152.060 ;
        RECT 1083.755 145.700 1084.140 151.485 ;
        RECT 1080.510 139.960 1080.845 141.310 ;
        RECT 1084.115 140.945 1084.540 145.220 ;
        RECT 1085.815 142.710 1086.115 149.750 ;
        RECT 1086.935 142.105 1087.235 149.035 ;
        RECT 1088.245 142.705 1088.545 149.055 ;
        RECT 1082.775 140.035 1083.155 140.415 ;
        RECT 1084.970 140.020 1085.350 140.400 ;
        RECT 1088.840 139.960 1089.130 149.740 ;
        RECT 1089.560 142.735 1089.855 149.560 ;
        RECT 1090.690 142.195 1090.990 149.005 ;
        RECT 1091.480 142.790 1091.790 152.830 ;
        RECT 1100.670 151.075 1101.050 151.455 ;
        RECT 1092.275 142.720 1092.575 149.550 ;
        RECT 1093.400 142.105 1093.700 149.045 ;
        RECT 1094.850 141.980 1095.130 145.015 ;
        RECT 1095.610 142.680 1095.890 149.040 ;
        RECT 1096.460 142.680 1096.760 149.500 ;
        RECT 1097.600 141.935 1097.900 149.090 ;
        RECT 1098.245 146.125 1098.625 146.505 ;
        RECT 1098.245 144.070 1098.625 144.450 ;
        RECT 1100.095 143.950 1100.410 148.275 ;
        RECT 1100.705 146.025 1100.985 147.555 ;
        RECT 1101.275 142.710 1101.575 149.750 ;
        RECT 1102.395 142.105 1102.695 149.035 ;
        RECT 1103.050 143.465 1103.350 147.525 ;
        RECT 1103.705 142.705 1104.005 149.055 ;
        RECT 1100.570 140.900 1100.950 141.280 ;
        RECT 1104.300 140.495 1104.590 149.740 ;
        RECT 1105.020 142.735 1105.315 149.560 ;
        RECT 1106.150 142.195 1106.450 149.005 ;
        RECT 1106.940 142.790 1107.250 151.525 ;
        RECT 1107.735 142.720 1108.035 149.550 ;
        RECT 1108.860 142.105 1109.160 149.045 ;
        RECT 1109.540 143.450 1109.820 147.540 ;
        RECT 1110.310 141.980 1110.590 145.015 ;
        RECT 1111.070 142.680 1111.350 149.040 ;
        RECT 1111.920 142.680 1112.220 149.500 ;
        RECT 1113.060 141.935 1113.360 149.090 ;
        RECT 1115.100 147.830 1115.475 156.030 ;
        RECT 1116.845 147.025 1117.145 158.020 ;
        RECT 1118.275 145.975 1118.655 156.230 ;
        RECT 1119.145 143.820 1119.580 157.395 ;
        RECT 1174.850 156.640 1175.365 166.690 ;
        RECT 1183.530 166.235 1183.910 166.615 ;
        RECT 1176.535 155.285 1177.120 166.065 ;
        RECT 1183.495 165.565 1183.875 165.945 ;
        RECT 1184.210 162.490 1184.510 169.530 ;
        RECT 1185.330 161.885 1185.630 168.815 ;
        RECT 1185.985 163.245 1186.285 167.305 ;
        RECT 1186.640 162.485 1186.940 168.835 ;
        RECT 1187.235 164.360 1187.555 169.520 ;
        RECT 1187.955 162.515 1188.250 169.340 ;
        RECT 1189.085 161.975 1189.385 168.785 ;
        RECT 1189.875 162.570 1190.185 168.760 ;
        RECT 1190.670 162.500 1190.970 169.330 ;
        RECT 1191.795 161.885 1192.095 168.825 ;
        RECT 1192.475 163.230 1192.755 167.320 ;
        RECT 1193.245 161.760 1193.525 164.795 ;
        RECT 1194.005 162.460 1194.310 168.820 ;
        RECT 1194.855 162.460 1195.155 169.280 ;
        RECT 1195.995 161.715 1196.295 168.870 ;
        RECT 1196.660 167.670 1197.040 168.050 ;
        RECT 1198.930 167.670 1199.310 168.075 ;
        RECT 1196.665 166.920 1197.045 167.300 ;
        RECT 1198.935 166.920 1199.315 167.325 ;
        RECT 1196.665 165.905 1197.045 166.285 ;
        RECT 1198.450 164.485 1198.770 166.615 ;
        RECT 1196.880 161.195 1197.260 164.215 ;
        RECT 1199.060 163.645 1199.340 166.050 ;
        RECT 1199.670 162.490 1199.970 169.530 ;
        RECT 1200.790 161.885 1201.090 168.815 ;
        RECT 1201.445 163.245 1201.745 167.305 ;
        RECT 1202.100 162.485 1202.400 168.835 ;
        RECT 1202.695 164.360 1203.020 169.520 ;
        RECT 1203.415 162.515 1203.710 169.340 ;
        RECT 1204.545 161.975 1204.845 168.785 ;
        RECT 1205.335 162.570 1205.645 168.760 ;
        RECT 1206.130 162.500 1206.430 169.330 ;
        RECT 1207.255 161.885 1207.555 168.825 ;
        RECT 1207.935 163.230 1208.215 167.320 ;
        RECT 1208.705 161.760 1208.985 164.795 ;
        RECT 1209.465 162.460 1209.785 168.820 ;
        RECT 1210.315 162.460 1210.615 169.280 ;
        RECT 1211.455 161.715 1211.755 168.870 ;
        RECT 1212.395 167.670 1212.755 169.500 ;
        RECT 1212.090 163.860 1212.470 164.240 ;
        RECT 1212.795 159.745 1213.155 166.305 ;
        RECT 1213.935 164.495 1214.260 166.360 ;
        RECT 1214.575 166.150 1214.990 169.500 ;
        RECT 1214.600 161.150 1215.060 165.835 ;
        RECT 1215.385 163.695 1215.835 172.515 ;
        RECT 1216.245 161.320 1216.600 171.625 ;
        RECT 1216.910 166.925 1217.255 167.980 ;
        RECT 1217.570 165.520 1218.000 168.510 ;
        RECT 1215.315 159.805 1215.695 160.185 ;
        RECT 1218.205 159.825 1218.585 161.200 ;
        RECT 1218.975 160.645 1219.290 171.695 ;
        RECT 1219.990 170.390 1220.280 172.450 ;
        RECT 1222.775 170.990 1223.250 174.040 ;
        RECT 1227.730 170.900 1228.140 173.995 ;
        RECT 1226.770 169.240 1227.080 169.270 ;
        RECT 1219.910 162.535 1220.235 164.905 ;
        RECT 1221.560 164.580 1221.960 168.545 ;
        RECT 1220.645 158.795 1220.990 161.255 ;
        RECT 1222.280 160.475 1222.605 163.240 ;
        RECT 1223.265 162.510 1223.670 165.840 ;
        RECT 1226.770 163.140 1227.085 169.240 ;
        RECT 1227.915 159.535 1228.285 168.635 ;
        RECT 1228.860 160.600 1229.150 172.435 ;
        RECT 1232.310 170.875 1232.720 173.970 ;
        RECT 1236.765 170.330 1237.075 172.845 ;
        RECT 1229.755 163.095 1230.085 169.290 ;
        RECT 1232.675 162.565 1233.115 165.840 ;
        RECT 1235.055 164.580 1235.580 168.520 ;
        RECT 1234.215 160.475 1234.540 163.240 ;
        RECT 1236.730 162.570 1237.145 164.960 ;
        RECT 1237.760 161.130 1238.075 171.815 ;
        RECT 1239.090 165.520 1239.575 168.530 ;
        RECT 1240.270 161.145 1240.600 171.840 ;
        RECT 1238.460 159.740 1238.795 161.090 ;
        RECT 1150.035 140.980 1150.350 152.030 ;
        RECT 1153.870 151.325 1154.270 154.375 ;
        RECT 1158.790 151.235 1159.200 154.330 ;
        RECT 1163.370 151.210 1163.780 154.305 ;
        RECT 1151.705 139.130 1152.050 141.590 ;
        RECT 1168.820 141.465 1169.135 152.150 ;
        RECT 1174.005 144.255 1174.455 148.415 ;
        RECT 1175.705 147.235 1176.230 147.675 ;
        RECT 987.300 128.270 987.680 128.650 ;
        RECT 987.290 127.520 987.670 127.900 ;
        RECT 987.335 126.835 987.715 127.215 ;
        RECT 987.300 126.165 987.680 126.545 ;
        RECT 988.015 123.090 988.315 130.130 ;
        RECT 989.135 122.485 989.435 129.415 ;
        RECT 989.790 123.845 990.090 127.905 ;
        RECT 990.445 123.085 990.745 129.435 ;
        RECT 991.040 124.960 991.360 130.120 ;
        RECT 991.760 123.115 992.055 129.940 ;
        RECT 992.890 122.575 993.190 129.385 ;
        RECT 993.680 123.170 993.990 129.360 ;
        RECT 994.475 123.100 994.775 129.930 ;
        RECT 995.600 122.485 995.900 129.425 ;
        RECT 996.280 123.830 996.560 127.920 ;
        RECT 997.050 122.360 997.330 125.395 ;
        RECT 997.810 123.060 998.115 129.420 ;
        RECT 998.660 123.060 998.960 129.880 ;
        RECT 999.800 122.315 1000.100 129.470 ;
        RECT 1000.465 128.270 1000.845 128.650 ;
        RECT 1002.735 128.270 1003.115 128.675 ;
        RECT 1000.470 127.520 1000.850 127.900 ;
        RECT 1002.740 127.520 1003.120 127.925 ;
        RECT 1000.470 126.505 1000.850 126.885 ;
        RECT 1002.255 125.085 1002.575 127.215 ;
        RECT 1000.685 121.795 1001.065 124.815 ;
        RECT 1002.865 124.245 1003.145 126.650 ;
        RECT 1003.475 123.090 1003.775 130.130 ;
        RECT 1004.595 122.485 1004.895 129.415 ;
        RECT 1005.250 123.845 1005.550 127.905 ;
        RECT 1005.905 123.085 1006.205 129.435 ;
        RECT 1006.500 124.960 1006.825 130.120 ;
        RECT 1007.220 123.115 1007.515 129.940 ;
        RECT 1008.350 122.575 1008.650 129.385 ;
        RECT 1009.140 123.170 1009.450 129.360 ;
        RECT 1009.935 123.100 1010.235 129.930 ;
        RECT 1011.060 122.485 1011.360 129.425 ;
        RECT 1011.740 123.830 1012.020 127.920 ;
        RECT 1012.510 122.360 1012.790 125.395 ;
        RECT 1013.270 123.060 1013.590 129.420 ;
        RECT 1014.120 123.060 1014.420 129.880 ;
        RECT 1015.260 122.315 1015.560 129.470 ;
        RECT 1016.200 128.270 1016.560 130.100 ;
        RECT 1015.895 124.460 1016.275 124.840 ;
        RECT 1016.600 120.345 1016.960 126.905 ;
        RECT 1017.740 125.095 1018.065 126.960 ;
        RECT 1018.380 126.750 1018.795 130.100 ;
        RECT 1018.405 121.750 1018.865 126.435 ;
        RECT 1019.190 124.295 1019.640 133.115 ;
        RECT 1020.050 121.920 1020.405 132.225 ;
        RECT 1020.715 127.525 1021.060 128.580 ;
        RECT 1021.375 126.120 1021.805 129.110 ;
        RECT 1019.120 120.405 1019.500 120.785 ;
        RECT 1022.010 120.425 1022.390 121.800 ;
        RECT 1022.780 121.245 1023.095 132.295 ;
        RECT 1023.795 130.990 1024.085 133.050 ;
        RECT 1026.580 131.590 1027.055 134.640 ;
        RECT 1031.535 131.500 1031.945 134.595 ;
        RECT 1030.575 129.840 1030.885 129.870 ;
        RECT 1023.715 123.135 1024.040 125.505 ;
        RECT 1025.365 125.180 1025.765 129.145 ;
        RECT 1024.450 119.395 1024.795 121.855 ;
        RECT 1026.085 121.075 1026.410 123.840 ;
        RECT 1027.070 123.110 1027.475 126.440 ;
        RECT 1030.575 123.740 1030.890 129.840 ;
        RECT 1031.720 120.135 1032.090 129.235 ;
        RECT 1032.665 121.200 1032.955 133.035 ;
        RECT 1036.115 131.475 1036.525 134.570 ;
        RECT 1040.570 130.930 1040.880 133.445 ;
        RECT 1033.560 123.695 1033.890 129.890 ;
        RECT 1036.480 123.165 1036.920 126.440 ;
        RECT 1038.860 125.180 1039.385 129.120 ;
        RECT 1038.020 121.075 1038.345 123.840 ;
        RECT 1040.535 123.170 1040.950 125.560 ;
        RECT 1041.565 121.730 1041.880 132.415 ;
        RECT 1042.895 126.120 1043.380 129.130 ;
        RECT 1044.075 121.745 1044.405 132.440 ;
        RECT 1042.265 120.340 1042.600 121.690 ;
        RECT 953.700 101.400 954.015 112.450 ;
        RECT 957.535 111.745 957.935 114.795 ;
        RECT 962.455 111.655 962.865 114.750 ;
        RECT 967.035 111.630 967.445 114.725 ;
        RECT 955.370 99.550 955.715 102.010 ;
        RECT 972.485 101.885 972.800 112.570 ;
        RECT 977.670 104.675 978.120 108.835 ;
        RECT 979.370 107.655 979.895 108.095 ;
        RECT 790.635 88.720 791.015 89.100 ;
        RECT 790.625 87.970 791.005 88.350 ;
        RECT 790.670 87.285 791.050 87.665 ;
        RECT 790.635 86.615 791.015 86.995 ;
        RECT 791.350 83.540 791.650 90.580 ;
        RECT 792.470 82.935 792.770 89.865 ;
        RECT 793.125 84.295 793.425 88.355 ;
        RECT 793.780 83.535 794.080 89.885 ;
        RECT 794.375 85.410 794.695 90.570 ;
        RECT 795.095 83.565 795.390 90.390 ;
        RECT 796.225 83.025 796.525 89.835 ;
        RECT 797.015 83.620 797.325 89.810 ;
        RECT 797.810 83.550 798.110 90.380 ;
        RECT 798.935 82.935 799.235 89.875 ;
        RECT 799.615 84.280 799.895 88.370 ;
        RECT 800.385 82.810 800.665 85.845 ;
        RECT 801.145 83.510 801.450 89.870 ;
        RECT 801.995 83.510 802.295 90.330 ;
        RECT 803.135 82.765 803.435 89.920 ;
        RECT 803.800 88.720 804.180 89.100 ;
        RECT 806.070 88.720 806.450 89.125 ;
        RECT 803.805 87.970 804.185 88.350 ;
        RECT 806.075 87.970 806.455 88.375 ;
        RECT 803.805 86.955 804.185 87.335 ;
        RECT 805.590 85.535 805.910 87.665 ;
        RECT 804.020 82.245 804.400 85.265 ;
        RECT 806.200 84.695 806.480 87.100 ;
        RECT 806.810 83.540 807.110 90.580 ;
        RECT 807.930 82.935 808.230 89.865 ;
        RECT 808.585 84.295 808.885 88.355 ;
        RECT 809.240 83.535 809.540 89.885 ;
        RECT 809.835 85.410 810.160 90.570 ;
        RECT 810.555 83.565 810.850 90.390 ;
        RECT 811.685 83.025 811.985 89.835 ;
        RECT 812.475 83.620 812.785 89.810 ;
        RECT 813.270 83.550 813.570 90.380 ;
        RECT 814.395 82.935 814.695 89.875 ;
        RECT 815.075 84.280 815.355 88.370 ;
        RECT 815.845 82.810 816.125 85.845 ;
        RECT 816.605 83.510 816.925 89.870 ;
        RECT 817.455 83.510 817.755 90.330 ;
        RECT 818.595 82.765 818.895 89.920 ;
        RECT 819.535 88.720 819.895 90.550 ;
        RECT 819.230 84.910 819.610 85.290 ;
        RECT 819.935 80.795 820.295 87.355 ;
        RECT 821.075 85.545 821.400 87.410 ;
        RECT 821.715 87.200 822.130 90.550 ;
        RECT 821.740 82.200 822.200 86.885 ;
        RECT 822.525 84.745 822.975 93.565 ;
        RECT 823.385 82.370 823.740 92.675 ;
        RECT 824.050 87.975 824.395 89.030 ;
        RECT 824.710 86.570 825.140 89.560 ;
        RECT 822.455 80.855 822.835 81.235 ;
        RECT 825.345 80.875 825.725 82.250 ;
        RECT 826.115 81.695 826.430 92.745 ;
        RECT 827.130 91.440 827.420 93.500 ;
        RECT 829.915 92.040 830.390 95.090 ;
        RECT 834.870 91.950 835.280 95.045 ;
        RECT 833.910 90.290 834.220 90.320 ;
        RECT 827.050 83.585 827.375 85.955 ;
        RECT 828.700 85.630 829.100 89.595 ;
        RECT 827.785 79.845 828.130 82.305 ;
        RECT 829.420 81.525 829.745 84.290 ;
        RECT 830.405 83.560 830.810 86.890 ;
        RECT 833.910 84.190 834.225 90.290 ;
        RECT 835.055 80.585 835.425 89.685 ;
        RECT 836.000 81.650 836.290 93.485 ;
        RECT 839.450 91.925 839.860 95.020 ;
        RECT 843.905 91.380 844.215 93.895 ;
        RECT 836.895 84.145 837.225 90.340 ;
        RECT 839.815 83.615 840.255 86.890 ;
        RECT 842.195 85.630 842.720 89.570 ;
        RECT 841.355 81.525 841.680 84.290 ;
        RECT 843.870 83.620 844.285 86.010 ;
        RECT 844.900 82.180 845.215 92.865 ;
        RECT 846.230 86.570 846.715 89.580 ;
        RECT 847.410 82.195 847.740 92.890 ;
        RECT 845.600 80.790 845.935 82.140 ;
        RECT 757.275 61.860 757.590 72.910 ;
        RECT 761.110 72.205 761.510 75.255 ;
        RECT 766.030 72.115 766.440 75.210 ;
        RECT 770.610 72.090 771.020 75.185 ;
        RECT 758.945 60.010 759.290 62.470 ;
        RECT 776.060 62.345 776.375 73.030 ;
        RECT 781.245 65.135 781.695 69.295 ;
        RECT 782.945 68.115 783.470 68.555 ;
        RECT 594.375 49.150 594.755 49.530 ;
        RECT 594.365 48.400 594.745 48.780 ;
        RECT 594.410 47.715 594.790 48.095 ;
        RECT 594.375 47.045 594.755 47.425 ;
        RECT 595.090 43.970 595.390 51.010 ;
        RECT 596.210 43.365 596.510 50.295 ;
        RECT 596.865 44.725 597.165 48.785 ;
        RECT 597.520 43.965 597.820 50.315 ;
        RECT 598.115 45.840 598.435 51.000 ;
        RECT 598.835 43.995 599.130 50.820 ;
        RECT 599.965 43.455 600.265 50.265 ;
        RECT 600.755 44.050 601.065 50.240 ;
        RECT 601.550 43.980 601.850 50.810 ;
        RECT 602.675 43.365 602.975 50.305 ;
        RECT 603.355 44.710 603.635 48.800 ;
        RECT 604.125 43.240 604.405 46.275 ;
        RECT 604.885 43.940 605.190 50.300 ;
        RECT 605.735 43.940 606.035 50.760 ;
        RECT 606.875 43.195 607.175 50.350 ;
        RECT 607.540 49.150 607.920 49.530 ;
        RECT 609.810 49.150 610.190 49.555 ;
        RECT 607.545 48.400 607.925 48.780 ;
        RECT 609.815 48.400 610.195 48.805 ;
        RECT 607.545 47.385 607.925 47.765 ;
        RECT 609.330 45.965 609.650 48.095 ;
        RECT 607.760 42.675 608.140 45.695 ;
        RECT 609.940 45.125 610.220 47.530 ;
        RECT 610.550 43.970 610.850 51.010 ;
        RECT 611.670 43.365 611.970 50.295 ;
        RECT 612.325 44.725 612.625 48.785 ;
        RECT 612.980 43.965 613.280 50.315 ;
        RECT 613.575 45.840 613.900 51.000 ;
        RECT 614.295 43.995 614.590 50.820 ;
        RECT 615.425 43.455 615.725 50.265 ;
        RECT 616.215 44.050 616.525 50.240 ;
        RECT 617.010 43.980 617.310 50.810 ;
        RECT 618.135 43.365 618.435 50.305 ;
        RECT 618.815 44.710 619.095 48.800 ;
        RECT 619.585 43.240 619.865 46.275 ;
        RECT 620.345 43.940 620.665 50.300 ;
        RECT 621.195 43.940 621.495 50.760 ;
        RECT 622.335 43.195 622.635 50.350 ;
        RECT 623.275 49.150 623.635 50.980 ;
        RECT 622.970 45.340 623.350 45.720 ;
        RECT 623.675 41.225 624.035 47.785 ;
        RECT 624.815 45.975 625.140 47.840 ;
        RECT 625.455 47.630 625.870 50.980 ;
        RECT 625.480 42.630 625.940 47.315 ;
        RECT 626.265 45.175 626.715 53.995 ;
        RECT 627.125 42.800 627.480 53.105 ;
        RECT 627.790 48.405 628.135 49.460 ;
        RECT 628.450 47.000 628.880 49.990 ;
        RECT 626.195 41.285 626.575 41.665 ;
        RECT 629.085 41.305 629.465 42.680 ;
        RECT 629.855 42.125 630.170 53.175 ;
        RECT 630.870 51.870 631.160 53.930 ;
        RECT 633.655 52.470 634.130 55.520 ;
        RECT 638.610 52.380 639.020 55.475 ;
        RECT 637.650 50.720 637.960 50.750 ;
        RECT 630.790 44.015 631.115 46.385 ;
        RECT 632.440 46.060 632.840 50.025 ;
        RECT 631.525 40.275 631.870 42.735 ;
        RECT 633.160 41.955 633.485 44.720 ;
        RECT 634.145 43.990 634.550 47.320 ;
        RECT 637.650 44.620 637.965 50.720 ;
        RECT 638.795 41.015 639.165 50.115 ;
        RECT 639.740 42.080 640.030 53.915 ;
        RECT 643.190 52.355 643.600 55.450 ;
        RECT 647.645 51.810 647.955 54.325 ;
        RECT 640.635 44.575 640.965 50.770 ;
        RECT 643.555 44.045 643.995 47.320 ;
        RECT 645.935 46.060 646.460 50.000 ;
        RECT 645.095 41.955 645.420 44.720 ;
        RECT 647.610 44.050 648.025 46.440 ;
        RECT 648.640 42.610 648.955 53.295 ;
        RECT 649.970 47.000 650.455 50.010 ;
        RECT 651.150 42.625 651.480 53.320 ;
        RECT 649.340 41.220 649.675 42.570 ;
        RECT 560.955 22.405 561.270 33.455 ;
        RECT 564.790 32.750 565.190 35.800 ;
        RECT 569.710 32.660 570.120 35.755 ;
        RECT 574.290 32.635 574.700 35.730 ;
        RECT 562.625 20.555 562.970 23.015 ;
        RECT 579.740 22.890 580.055 33.575 ;
        RECT 584.975 25.605 585.425 29.765 ;
        RECT 586.675 28.585 587.200 29.025 ;
        RECT 469.440 3.790 469.740 10.720 ;
        RECT 470.095 5.150 470.395 9.210 ;
        RECT 470.750 4.390 471.050 10.740 ;
        RECT 472.065 4.420 472.360 11.245 ;
        RECT 475.905 3.790 476.205 10.730 ;
        RECT 476.585 5.135 476.865 9.225 ;
        RECT 478.115 4.365 478.420 10.725 ;
        RECT 478.965 4.365 479.265 11.185 ;
        RECT 480.695 7.805 481.075 8.185 ;
        RECT 480.705 5.760 481.085 6.140 ;
        RECT 585.775 5.445 586.290 27.690 ;
        RECT 587.460 7.660 588.045 28.415 ;
        RECT 589.110 25.220 589.465 39.160 ;
        RECT 652.455 38.530 652.905 48.795 ;
        RECT 590.735 26.010 591.095 37.560 ;
        RECT 653.620 36.990 654.105 45.875 ;
        RECT 660.560 36.265 660.965 48.310 ;
        RECT 662.635 38.165 663.025 49.590 ;
        RECT 665.795 42.005 666.150 53.090 ;
        RECT 669.540 51.730 669.830 53.790 ;
        RECT 672.310 52.330 672.810 55.380 ;
        RECT 677.280 52.240 677.690 55.335 ;
        RECT 676.320 50.580 676.630 50.610 ;
        RECT 667.120 46.860 667.590 49.850 ;
        RECT 669.470 43.875 669.785 46.245 ;
        RECT 671.090 45.920 671.510 49.885 ;
        RECT 667.755 41.165 668.135 42.540 ;
        RECT 670.195 40.135 670.540 42.595 ;
        RECT 671.830 41.815 672.155 44.580 ;
        RECT 672.815 43.850 673.220 47.180 ;
        RECT 676.320 44.480 676.635 50.580 ;
        RECT 677.465 40.875 677.835 49.975 ;
        RECT 678.410 41.940 678.700 53.775 ;
        RECT 681.860 52.215 682.270 55.310 ;
        RECT 686.315 51.670 686.625 54.185 ;
        RECT 690.565 53.370 690.945 53.750 ;
        RECT 692.695 53.370 693.075 53.750 ;
        RECT 679.305 44.435 679.635 50.630 ;
        RECT 682.210 43.905 682.665 47.180 ;
        RECT 684.570 45.920 685.115 49.860 ;
        RECT 688.625 46.860 689.060 49.870 ;
        RECT 683.765 41.815 684.090 44.580 ;
        RECT 686.280 43.910 686.695 46.300 ;
        RECT 689.820 42.485 690.150 53.180 ;
        RECT 691.255 46.820 691.640 52.605 ;
        RECT 688.010 41.080 688.345 42.430 ;
        RECT 691.615 42.065 692.040 46.340 ;
        RECT 693.315 43.830 693.615 50.870 ;
        RECT 694.435 43.225 694.735 50.155 ;
        RECT 695.745 43.825 696.045 50.175 ;
        RECT 690.275 41.155 690.655 41.535 ;
        RECT 692.470 41.140 692.850 41.520 ;
        RECT 696.340 41.080 696.630 50.860 ;
        RECT 697.060 43.855 697.355 50.680 ;
        RECT 698.190 43.315 698.490 50.125 ;
        RECT 698.980 43.910 699.290 53.950 ;
        RECT 708.170 52.195 708.550 52.575 ;
        RECT 699.775 43.840 700.075 50.670 ;
        RECT 700.900 43.225 701.200 50.165 ;
        RECT 702.350 43.100 702.630 46.135 ;
        RECT 703.110 43.800 703.390 50.160 ;
        RECT 703.960 43.800 704.260 50.620 ;
        RECT 705.100 43.055 705.400 50.210 ;
        RECT 705.745 47.245 706.125 47.625 ;
        RECT 705.745 45.190 706.125 45.570 ;
        RECT 707.595 45.070 707.910 49.395 ;
        RECT 708.205 47.145 708.485 48.675 ;
        RECT 708.775 43.830 709.075 50.870 ;
        RECT 709.895 43.225 710.195 50.155 ;
        RECT 710.550 44.585 710.850 48.645 ;
        RECT 711.205 43.825 711.505 50.175 ;
        RECT 708.070 42.020 708.450 42.400 ;
        RECT 711.800 41.615 712.090 50.860 ;
        RECT 712.520 43.855 712.815 50.680 ;
        RECT 713.650 43.315 713.950 50.125 ;
        RECT 714.440 43.910 714.750 52.645 ;
        RECT 715.235 43.840 715.535 50.670 ;
        RECT 716.360 43.225 716.660 50.165 ;
        RECT 717.040 44.570 717.320 48.660 ;
        RECT 717.810 43.100 718.090 46.135 ;
        RECT 718.570 43.800 718.850 50.160 ;
        RECT 719.420 43.800 719.720 50.620 ;
        RECT 720.560 43.055 720.860 50.210 ;
        RECT 722.900 48.825 723.275 57.025 ;
        RECT 724.645 48.020 724.945 59.015 ;
        RECT 725.565 47.105 725.945 57.360 ;
        RECT 726.435 44.950 726.870 58.525 ;
        RECT 782.145 57.685 782.660 67.985 ;
        RECT 783.830 56.580 784.415 67.360 ;
        RECT 785.355 64.825 785.710 78.745 ;
        RECT 848.700 78.115 849.150 88.380 ;
        RECT 786.980 65.730 787.340 77.145 ;
        RECT 849.865 76.575 850.350 85.460 ;
        RECT 856.530 76.310 856.935 87.840 ;
        RECT 858.605 78.210 858.995 89.310 ;
        RECT 862.030 81.690 862.385 92.775 ;
        RECT 865.775 91.415 866.065 93.475 ;
        RECT 868.545 92.015 869.045 95.065 ;
        RECT 873.515 91.925 873.925 95.020 ;
        RECT 872.555 90.265 872.865 90.295 ;
        RECT 863.355 86.545 863.825 89.535 ;
        RECT 865.705 83.560 866.020 85.930 ;
        RECT 867.325 85.605 867.745 89.570 ;
        RECT 863.990 80.850 864.370 82.225 ;
        RECT 866.430 79.820 866.775 82.280 ;
        RECT 868.065 81.500 868.390 84.265 ;
        RECT 869.050 83.535 869.455 86.865 ;
        RECT 872.555 84.165 872.870 90.265 ;
        RECT 873.700 80.560 874.070 89.660 ;
        RECT 874.645 81.625 874.935 93.460 ;
        RECT 878.095 91.900 878.505 94.995 ;
        RECT 882.550 91.355 882.860 93.870 ;
        RECT 886.800 93.055 887.180 93.435 ;
        RECT 888.930 93.055 889.310 93.435 ;
        RECT 875.540 84.120 875.870 90.315 ;
        RECT 878.445 83.590 878.900 86.865 ;
        RECT 880.805 85.605 881.350 89.545 ;
        RECT 884.860 86.545 885.295 89.555 ;
        RECT 880.000 81.500 880.325 84.265 ;
        RECT 882.515 83.595 882.930 85.985 ;
        RECT 886.055 82.170 886.385 92.865 ;
        RECT 887.490 86.505 887.875 92.290 ;
        RECT 884.245 80.765 884.580 82.115 ;
        RECT 887.850 81.750 888.275 86.025 ;
        RECT 889.550 83.515 889.850 90.555 ;
        RECT 890.670 82.910 890.970 89.840 ;
        RECT 891.980 83.510 892.280 89.860 ;
        RECT 886.510 80.840 886.890 81.220 ;
        RECT 888.705 80.825 889.085 81.205 ;
        RECT 892.575 80.765 892.865 90.545 ;
        RECT 893.295 83.540 893.590 90.365 ;
        RECT 894.425 83.000 894.725 89.810 ;
        RECT 895.215 83.595 895.525 93.635 ;
        RECT 904.405 91.880 904.785 92.260 ;
        RECT 896.010 83.525 896.310 90.355 ;
        RECT 897.135 82.910 897.435 89.850 ;
        RECT 898.585 82.785 898.865 85.820 ;
        RECT 899.345 83.485 899.625 89.845 ;
        RECT 900.195 83.485 900.495 90.305 ;
        RECT 901.335 82.740 901.635 89.895 ;
        RECT 901.980 86.930 902.360 87.310 ;
        RECT 901.980 84.875 902.360 85.255 ;
        RECT 903.830 84.755 904.145 89.080 ;
        RECT 904.440 86.830 904.720 88.360 ;
        RECT 905.010 83.515 905.310 90.555 ;
        RECT 906.130 82.910 906.430 89.840 ;
        RECT 906.785 84.270 907.085 88.330 ;
        RECT 907.440 83.510 907.740 89.860 ;
        RECT 904.305 81.705 904.685 82.085 ;
        RECT 908.035 81.300 908.325 90.545 ;
        RECT 908.755 83.540 909.050 90.365 ;
        RECT 909.885 83.000 910.185 89.810 ;
        RECT 910.675 83.595 910.985 92.330 ;
        RECT 911.470 83.525 911.770 90.355 ;
        RECT 912.595 82.910 912.895 89.850 ;
        RECT 913.275 84.255 913.555 88.345 ;
        RECT 914.045 82.785 914.325 85.820 ;
        RECT 914.805 83.485 915.085 89.845 ;
        RECT 915.655 83.485 915.955 90.305 ;
        RECT 916.795 82.740 917.095 89.895 ;
        RECT 919.080 88.600 919.455 96.885 ;
        RECT 920.825 87.880 921.125 98.875 ;
        RECT 921.950 86.775 922.330 97.030 ;
        RECT 922.820 84.620 923.255 98.195 ;
        RECT 978.525 97.395 979.040 107.445 ;
        RECT 980.210 96.040 980.795 106.820 ;
        RECT 982.045 104.375 982.400 118.165 ;
        RECT 1045.390 117.535 1045.840 128.035 ;
        RECT 983.670 105.230 984.030 116.565 ;
        RECT 1046.555 115.995 1047.040 125.235 ;
        RECT 1052.970 115.750 1053.375 127.280 ;
        RECT 1055.045 117.650 1055.435 128.750 ;
        RECT 1058.450 121.240 1058.805 132.325 ;
        RECT 1062.195 130.965 1062.485 133.025 ;
        RECT 1064.965 131.565 1065.465 134.615 ;
        RECT 1069.935 131.475 1070.345 134.570 ;
        RECT 1068.975 129.815 1069.285 129.845 ;
        RECT 1059.775 126.095 1060.245 129.085 ;
        RECT 1062.125 123.110 1062.440 125.480 ;
        RECT 1063.745 125.155 1064.165 129.120 ;
        RECT 1060.410 120.400 1060.790 121.775 ;
        RECT 1062.850 119.370 1063.195 121.830 ;
        RECT 1064.485 121.050 1064.810 123.815 ;
        RECT 1065.470 123.085 1065.875 126.415 ;
        RECT 1068.975 123.715 1069.290 129.815 ;
        RECT 1070.120 120.110 1070.490 129.210 ;
        RECT 1071.065 121.175 1071.355 133.010 ;
        RECT 1074.515 131.450 1074.925 134.545 ;
        RECT 1078.970 130.905 1079.280 133.420 ;
        RECT 1083.220 132.605 1083.600 132.985 ;
        RECT 1085.350 132.605 1085.730 132.985 ;
        RECT 1071.960 123.670 1072.290 129.865 ;
        RECT 1074.865 123.140 1075.320 126.415 ;
        RECT 1077.225 125.155 1077.770 129.095 ;
        RECT 1081.280 126.095 1081.715 129.105 ;
        RECT 1076.420 121.050 1076.745 123.815 ;
        RECT 1078.935 123.145 1079.350 125.535 ;
        RECT 1082.475 121.720 1082.805 132.415 ;
        RECT 1083.910 126.055 1084.295 131.840 ;
        RECT 1080.665 120.315 1081.000 121.665 ;
        RECT 1084.270 121.300 1084.695 125.575 ;
        RECT 1085.970 123.065 1086.270 130.105 ;
        RECT 1087.090 122.460 1087.390 129.390 ;
        RECT 1088.400 123.060 1088.700 129.410 ;
        RECT 1082.930 120.390 1083.310 120.770 ;
        RECT 1085.125 120.375 1085.505 120.755 ;
        RECT 1088.995 120.315 1089.285 130.095 ;
        RECT 1089.715 123.090 1090.010 129.915 ;
        RECT 1090.845 122.550 1091.145 129.360 ;
        RECT 1091.635 123.145 1091.945 133.185 ;
        RECT 1100.825 131.430 1101.205 131.810 ;
        RECT 1092.430 123.075 1092.730 129.905 ;
        RECT 1093.555 122.460 1093.855 129.400 ;
        RECT 1095.005 122.335 1095.285 125.370 ;
        RECT 1095.765 123.035 1096.045 129.395 ;
        RECT 1096.615 123.035 1096.915 129.855 ;
        RECT 1097.755 122.290 1098.055 129.445 ;
        RECT 1098.400 126.480 1098.780 126.860 ;
        RECT 1098.400 124.425 1098.780 124.805 ;
        RECT 1100.250 124.305 1100.565 128.630 ;
        RECT 1100.860 126.380 1101.140 127.910 ;
        RECT 1101.430 123.065 1101.730 130.105 ;
        RECT 1102.550 122.460 1102.850 129.390 ;
        RECT 1103.205 123.820 1103.505 127.880 ;
        RECT 1103.860 123.060 1104.160 129.410 ;
        RECT 1100.725 121.255 1101.105 121.635 ;
        RECT 1104.455 120.850 1104.745 130.095 ;
        RECT 1105.175 123.090 1105.470 129.915 ;
        RECT 1106.305 122.550 1106.605 129.360 ;
        RECT 1107.095 123.145 1107.405 131.880 ;
        RECT 1107.890 123.075 1108.190 129.905 ;
        RECT 1109.015 122.460 1109.315 129.400 ;
        RECT 1109.695 123.805 1109.975 127.895 ;
        RECT 1110.465 122.335 1110.745 125.370 ;
        RECT 1111.225 123.035 1111.505 129.395 ;
        RECT 1112.075 123.035 1112.375 129.855 ;
        RECT 1113.215 122.290 1113.515 129.445 ;
        RECT 1115.400 128.080 1115.775 136.280 ;
        RECT 1117.145 127.275 1117.445 138.270 ;
        RECT 1118.275 126.330 1118.655 136.585 ;
        RECT 1119.145 124.175 1119.580 137.750 ;
        RECT 1174.850 136.950 1175.365 147.000 ;
        RECT 1176.535 135.595 1177.120 146.375 ;
        RECT 1178.175 143.915 1178.530 157.705 ;
        RECT 1241.520 157.075 1241.970 167.340 ;
        RECT 1179.800 144.770 1180.160 156.105 ;
        RECT 1242.685 155.535 1243.170 164.420 ;
        RECT 1248.990 155.160 1249.395 166.690 ;
        RECT 1251.065 157.060 1251.455 168.160 ;
        RECT 1254.835 160.610 1255.190 171.695 ;
        RECT 1256.160 165.465 1256.630 168.455 ;
        RECT 1256.795 159.770 1257.175 161.145 ;
        RECT 1257.565 160.590 1257.880 171.640 ;
        RECT 1258.580 170.335 1258.870 172.395 ;
        RECT 1261.350 170.935 1261.850 173.985 ;
        RECT 1266.320 170.845 1266.730 173.940 ;
        RECT 1265.360 169.185 1265.670 169.215 ;
        RECT 1258.510 162.480 1258.825 164.850 ;
        RECT 1260.130 164.525 1260.550 168.490 ;
        RECT 1259.235 158.740 1259.580 161.200 ;
        RECT 1260.870 160.420 1261.195 163.185 ;
        RECT 1261.855 162.455 1262.260 165.785 ;
        RECT 1265.360 163.085 1265.675 169.185 ;
        RECT 1266.505 159.480 1266.875 168.580 ;
        RECT 1267.450 160.545 1267.740 172.380 ;
        RECT 1270.900 170.820 1271.310 173.915 ;
        RECT 1275.355 170.275 1275.665 172.790 ;
        RECT 1279.605 171.975 1279.985 172.355 ;
        RECT 1281.735 171.975 1282.115 172.355 ;
        RECT 1268.345 163.040 1268.675 169.235 ;
        RECT 1271.250 162.510 1271.705 165.785 ;
        RECT 1273.610 164.525 1274.155 168.465 ;
        RECT 1272.805 160.420 1273.130 163.185 ;
        RECT 1275.320 162.515 1275.735 164.905 ;
        RECT 1276.350 161.075 1276.665 171.760 ;
        RECT 1277.665 165.465 1278.100 168.475 ;
        RECT 1278.860 161.090 1279.190 171.785 ;
        RECT 1279.540 166.835 1279.960 167.295 ;
        RECT 1280.295 165.425 1280.680 171.210 ;
        RECT 1281.040 166.830 1281.460 167.290 ;
        RECT 1279.675 163.945 1280.055 164.325 ;
        RECT 1277.050 159.685 1277.385 161.035 ;
        RECT 1280.655 160.670 1281.080 164.945 ;
        RECT 1281.740 163.920 1282.050 168.040 ;
        RECT 1282.355 162.435 1282.655 169.475 ;
        RECT 1283.475 161.830 1283.775 168.760 ;
        RECT 1284.130 163.190 1284.430 167.250 ;
        RECT 1284.785 162.430 1285.085 168.780 ;
        RECT 1279.315 159.760 1279.695 160.140 ;
        RECT 1281.510 159.745 1281.890 160.125 ;
        RECT 1285.380 159.685 1285.670 169.465 ;
        RECT 1286.100 162.460 1286.395 169.285 ;
        RECT 1287.230 161.920 1287.530 168.730 ;
        RECT 1288.020 162.515 1288.330 172.555 ;
        RECT 1288.815 162.445 1289.115 169.275 ;
        RECT 1289.940 161.830 1290.240 168.770 ;
        RECT 1290.620 163.175 1290.900 167.265 ;
        RECT 1291.390 161.705 1291.670 164.740 ;
        RECT 1292.150 162.405 1292.430 168.765 ;
        RECT 1293.000 162.405 1293.300 169.225 ;
        RECT 1294.140 161.660 1294.440 168.815 ;
        RECT 1294.810 167.615 1295.105 172.985 ;
        RECT 1295.385 166.785 1295.690 172.260 ;
        RECT 1297.210 170.800 1297.590 171.180 ;
        RECT 1294.785 165.850 1295.165 166.230 ;
        RECT 1294.785 163.795 1295.165 164.175 ;
        RECT 1296.635 163.675 1296.950 168.000 ;
        RECT 1297.245 165.750 1297.525 167.280 ;
        RECT 1297.815 162.435 1298.115 169.475 ;
        RECT 1299.590 163.190 1299.890 167.250 ;
        RECT 1297.110 160.625 1297.490 161.005 ;
        RECT 1300.840 160.220 1301.130 169.465 ;
        RECT 1302.690 161.920 1302.990 168.730 ;
        RECT 1303.480 162.515 1303.790 171.250 ;
        RECT 1304.275 162.445 1304.575 169.275 ;
        RECT 1306.080 163.175 1306.360 167.265 ;
        RECT 1306.850 161.705 1307.130 164.740 ;
        RECT 1309.600 161.660 1309.900 168.815 ;
        RECT 1183.450 147.980 1183.830 148.360 ;
        RECT 1183.440 147.230 1183.820 147.610 ;
        RECT 1183.485 146.545 1183.865 146.925 ;
        RECT 1183.450 145.875 1183.830 146.255 ;
        RECT 1184.165 142.800 1184.465 149.840 ;
        RECT 1185.285 142.195 1185.585 149.125 ;
        RECT 1185.940 143.555 1186.240 147.615 ;
        RECT 1186.595 142.795 1186.895 149.145 ;
        RECT 1187.190 144.670 1187.510 149.830 ;
        RECT 1187.910 142.825 1188.205 149.650 ;
        RECT 1189.040 142.285 1189.340 149.095 ;
        RECT 1189.830 142.880 1190.140 149.070 ;
        RECT 1190.625 142.810 1190.925 149.640 ;
        RECT 1191.750 142.195 1192.050 149.135 ;
        RECT 1192.430 143.540 1192.710 147.630 ;
        RECT 1193.200 142.070 1193.480 145.105 ;
        RECT 1193.960 142.770 1194.265 149.130 ;
        RECT 1194.810 142.770 1195.110 149.590 ;
        RECT 1195.950 142.025 1196.250 149.180 ;
        RECT 1196.615 147.980 1196.995 148.360 ;
        RECT 1198.885 147.980 1199.265 148.385 ;
        RECT 1196.620 147.230 1197.000 147.610 ;
        RECT 1198.890 147.230 1199.270 147.635 ;
        RECT 1196.620 146.215 1197.000 146.595 ;
        RECT 1198.405 144.795 1198.725 146.925 ;
        RECT 1196.835 141.505 1197.215 144.525 ;
        RECT 1199.015 143.955 1199.295 146.360 ;
        RECT 1199.625 142.800 1199.925 149.840 ;
        RECT 1200.745 142.195 1201.045 149.125 ;
        RECT 1201.400 143.555 1201.700 147.615 ;
        RECT 1202.055 142.795 1202.355 149.145 ;
        RECT 1202.650 144.670 1202.975 149.830 ;
        RECT 1203.370 142.825 1203.665 149.650 ;
        RECT 1204.500 142.285 1204.800 149.095 ;
        RECT 1205.290 142.880 1205.600 149.070 ;
        RECT 1206.085 142.810 1206.385 149.640 ;
        RECT 1207.210 142.195 1207.510 149.135 ;
        RECT 1207.890 143.540 1208.170 147.630 ;
        RECT 1208.660 142.070 1208.940 145.105 ;
        RECT 1209.420 142.770 1209.740 149.130 ;
        RECT 1210.270 142.770 1210.570 149.590 ;
        RECT 1211.410 142.025 1211.710 149.180 ;
        RECT 1212.350 147.980 1212.710 149.810 ;
        RECT 1212.045 144.170 1212.425 144.550 ;
        RECT 1212.750 140.055 1213.110 146.615 ;
        RECT 1213.890 144.805 1214.215 146.670 ;
        RECT 1214.530 146.460 1214.945 149.810 ;
        RECT 1214.555 141.460 1215.015 146.145 ;
        RECT 1215.340 144.005 1215.790 152.825 ;
        RECT 1216.200 141.630 1216.555 151.935 ;
        RECT 1216.865 147.235 1217.210 148.290 ;
        RECT 1217.525 145.830 1217.955 148.820 ;
        RECT 1215.270 140.115 1215.650 140.495 ;
        RECT 1218.160 140.135 1218.540 141.510 ;
        RECT 1218.930 140.955 1219.245 152.005 ;
        RECT 1219.945 150.700 1220.235 152.760 ;
        RECT 1222.730 151.300 1223.205 154.350 ;
        RECT 1227.685 151.210 1228.095 154.305 ;
        RECT 1226.725 149.550 1227.035 149.580 ;
        RECT 1219.865 142.845 1220.190 145.215 ;
        RECT 1221.515 144.890 1221.915 148.855 ;
        RECT 1220.600 139.105 1220.945 141.565 ;
        RECT 1222.235 140.785 1222.560 143.550 ;
        RECT 1223.220 142.820 1223.625 146.150 ;
        RECT 1226.725 143.450 1227.040 149.550 ;
        RECT 1227.870 139.845 1228.240 148.945 ;
        RECT 1228.815 140.910 1229.105 152.745 ;
        RECT 1232.265 151.185 1232.675 154.280 ;
        RECT 1236.720 150.640 1237.030 153.155 ;
        RECT 1229.710 143.405 1230.040 149.600 ;
        RECT 1232.630 142.875 1233.070 146.150 ;
        RECT 1235.010 144.890 1235.535 148.830 ;
        RECT 1234.170 140.785 1234.495 143.550 ;
        RECT 1236.685 142.880 1237.100 145.270 ;
        RECT 1237.715 141.440 1238.030 152.125 ;
        RECT 1239.045 145.830 1239.530 148.840 ;
        RECT 1240.225 141.455 1240.555 152.150 ;
        RECT 1238.415 140.050 1238.750 141.400 ;
        RECT 1150.095 121.175 1150.410 132.225 ;
        RECT 1153.930 131.520 1154.330 134.570 ;
        RECT 1158.850 131.430 1159.260 134.525 ;
        RECT 1163.430 131.405 1163.840 134.500 ;
        RECT 1151.765 119.325 1152.110 121.785 ;
        RECT 1168.880 121.660 1169.195 132.345 ;
        RECT 1174.065 124.450 1174.515 128.610 ;
        RECT 1175.765 127.430 1176.290 127.870 ;
        RECT 987.105 108.430 987.485 108.810 ;
        RECT 987.095 107.680 987.475 108.060 ;
        RECT 987.140 106.995 987.520 107.375 ;
        RECT 987.105 106.325 987.485 106.705 ;
        RECT 987.820 103.250 988.120 110.290 ;
        RECT 988.940 102.645 989.240 109.575 ;
        RECT 989.595 104.005 989.895 108.065 ;
        RECT 990.250 103.245 990.550 109.595 ;
        RECT 990.845 105.120 991.165 110.280 ;
        RECT 991.565 103.275 991.860 110.100 ;
        RECT 992.695 102.735 992.995 109.545 ;
        RECT 993.485 103.330 993.795 109.520 ;
        RECT 994.280 103.260 994.580 110.090 ;
        RECT 995.405 102.645 995.705 109.585 ;
        RECT 996.085 103.990 996.365 108.080 ;
        RECT 996.855 102.520 997.135 105.555 ;
        RECT 997.615 103.220 997.920 109.580 ;
        RECT 998.465 103.220 998.765 110.040 ;
        RECT 999.605 102.475 999.905 109.630 ;
        RECT 1000.270 108.430 1000.650 108.810 ;
        RECT 1002.540 108.430 1002.920 108.835 ;
        RECT 1000.275 107.680 1000.655 108.060 ;
        RECT 1002.545 107.680 1002.925 108.085 ;
        RECT 1000.275 106.665 1000.655 107.045 ;
        RECT 1002.060 105.245 1002.380 107.375 ;
        RECT 1000.490 101.955 1000.870 104.975 ;
        RECT 1002.670 104.405 1002.950 106.810 ;
        RECT 1003.280 103.250 1003.580 110.290 ;
        RECT 1004.400 102.645 1004.700 109.575 ;
        RECT 1005.055 104.005 1005.355 108.065 ;
        RECT 1005.710 103.245 1006.010 109.595 ;
        RECT 1006.305 105.120 1006.630 110.280 ;
        RECT 1007.025 103.275 1007.320 110.100 ;
        RECT 1008.155 102.735 1008.455 109.545 ;
        RECT 1008.945 103.330 1009.255 109.520 ;
        RECT 1009.740 103.260 1010.040 110.090 ;
        RECT 1010.865 102.645 1011.165 109.585 ;
        RECT 1011.545 103.990 1011.825 108.080 ;
        RECT 1012.315 102.520 1012.595 105.555 ;
        RECT 1013.075 103.220 1013.395 109.580 ;
        RECT 1013.925 103.220 1014.225 110.040 ;
        RECT 1015.065 102.475 1015.365 109.630 ;
        RECT 1016.005 108.430 1016.365 110.260 ;
        RECT 1015.700 104.620 1016.080 105.000 ;
        RECT 1016.405 100.505 1016.765 107.065 ;
        RECT 1017.545 105.255 1017.870 107.120 ;
        RECT 1018.185 106.910 1018.600 110.260 ;
        RECT 1018.210 101.910 1018.670 106.595 ;
        RECT 1018.995 104.455 1019.445 113.275 ;
        RECT 1019.855 102.080 1020.210 112.385 ;
        RECT 1020.520 107.685 1020.865 108.740 ;
        RECT 1021.180 106.280 1021.610 109.270 ;
        RECT 1018.925 100.565 1019.305 100.945 ;
        RECT 1021.815 100.585 1022.195 101.960 ;
        RECT 1022.585 101.405 1022.900 112.455 ;
        RECT 1023.600 111.150 1023.890 113.210 ;
        RECT 1026.385 111.750 1026.860 114.800 ;
        RECT 1031.340 111.660 1031.750 114.755 ;
        RECT 1030.380 110.000 1030.690 110.030 ;
        RECT 1023.520 103.295 1023.845 105.665 ;
        RECT 1025.170 105.340 1025.570 109.305 ;
        RECT 1024.255 99.555 1024.600 102.015 ;
        RECT 1025.890 101.235 1026.215 104.000 ;
        RECT 1026.875 103.270 1027.280 106.600 ;
        RECT 1030.380 103.900 1030.695 110.000 ;
        RECT 1031.525 100.295 1031.895 109.395 ;
        RECT 1032.470 101.360 1032.760 113.195 ;
        RECT 1035.920 111.635 1036.330 114.730 ;
        RECT 1040.375 111.090 1040.685 113.605 ;
        RECT 1033.365 103.855 1033.695 110.050 ;
        RECT 1036.285 103.325 1036.725 106.600 ;
        RECT 1038.665 105.340 1039.190 109.280 ;
        RECT 1037.825 101.235 1038.150 104.000 ;
        RECT 1040.340 103.330 1040.755 105.720 ;
        RECT 1041.370 101.890 1041.685 112.575 ;
        RECT 1042.700 106.280 1043.185 109.290 ;
        RECT 1043.880 101.905 1044.210 112.600 ;
        RECT 1042.070 100.500 1042.405 101.850 ;
        RECT 953.730 81.675 954.045 92.725 ;
        RECT 957.565 92.020 957.965 95.070 ;
        RECT 962.485 91.930 962.895 95.025 ;
        RECT 967.065 91.905 967.475 95.000 ;
        RECT 955.400 79.825 955.745 82.285 ;
        RECT 972.515 82.160 972.830 92.845 ;
        RECT 977.700 84.950 978.150 89.110 ;
        RECT 979.400 87.930 979.925 88.370 ;
        RECT 790.765 68.960 791.145 69.340 ;
        RECT 790.755 68.210 791.135 68.590 ;
        RECT 790.800 67.525 791.180 67.905 ;
        RECT 790.765 66.855 791.145 67.235 ;
        RECT 791.480 63.780 791.780 70.820 ;
        RECT 792.600 63.175 792.900 70.105 ;
        RECT 793.255 64.535 793.555 68.595 ;
        RECT 793.910 63.775 794.210 70.125 ;
        RECT 794.505 65.650 794.825 70.810 ;
        RECT 795.225 63.805 795.520 70.630 ;
        RECT 796.355 63.265 796.655 70.075 ;
        RECT 797.145 63.860 797.455 70.050 ;
        RECT 797.940 63.790 798.240 70.620 ;
        RECT 799.065 63.175 799.365 70.115 ;
        RECT 799.745 64.520 800.025 68.610 ;
        RECT 800.515 63.050 800.795 66.085 ;
        RECT 801.275 63.750 801.580 70.110 ;
        RECT 802.125 63.750 802.425 70.570 ;
        RECT 803.265 63.005 803.565 70.160 ;
        RECT 803.930 68.960 804.310 69.340 ;
        RECT 806.200 68.960 806.580 69.365 ;
        RECT 803.935 68.210 804.315 68.590 ;
        RECT 806.205 68.210 806.585 68.615 ;
        RECT 803.935 67.195 804.315 67.575 ;
        RECT 805.720 65.775 806.040 67.905 ;
        RECT 804.150 62.485 804.530 65.505 ;
        RECT 806.330 64.935 806.610 67.340 ;
        RECT 806.940 63.780 807.240 70.820 ;
        RECT 808.060 63.175 808.360 70.105 ;
        RECT 808.715 64.535 809.015 68.595 ;
        RECT 809.370 63.775 809.670 70.125 ;
        RECT 809.965 65.650 810.290 70.810 ;
        RECT 810.685 63.805 810.980 70.630 ;
        RECT 811.815 63.265 812.115 70.075 ;
        RECT 812.605 63.860 812.915 70.050 ;
        RECT 813.400 63.790 813.700 70.620 ;
        RECT 814.525 63.175 814.825 70.115 ;
        RECT 815.205 64.520 815.485 68.610 ;
        RECT 815.975 63.050 816.255 66.085 ;
        RECT 816.735 63.750 817.055 70.110 ;
        RECT 817.585 63.750 817.885 70.570 ;
        RECT 818.725 63.005 819.025 70.160 ;
        RECT 819.665 68.960 820.025 70.790 ;
        RECT 819.360 65.150 819.740 65.530 ;
        RECT 820.065 61.035 820.425 67.595 ;
        RECT 821.205 65.785 821.530 67.650 ;
        RECT 821.845 67.440 822.260 70.790 ;
        RECT 821.870 62.440 822.330 67.125 ;
        RECT 822.655 64.985 823.105 73.805 ;
        RECT 823.515 62.610 823.870 72.915 ;
        RECT 824.180 68.215 824.525 69.270 ;
        RECT 824.840 66.810 825.270 69.800 ;
        RECT 822.585 61.095 822.965 61.475 ;
        RECT 825.475 61.115 825.855 62.490 ;
        RECT 826.245 61.935 826.560 72.985 ;
        RECT 827.260 71.680 827.550 73.740 ;
        RECT 830.045 72.280 830.520 75.330 ;
        RECT 835.000 72.190 835.410 75.285 ;
        RECT 834.040 70.530 834.350 70.560 ;
        RECT 827.180 63.825 827.505 66.195 ;
        RECT 828.830 65.870 829.230 69.835 ;
        RECT 827.915 60.085 828.260 62.545 ;
        RECT 829.550 61.765 829.875 64.530 ;
        RECT 830.535 63.800 830.940 67.130 ;
        RECT 834.040 64.430 834.355 70.530 ;
        RECT 835.185 60.825 835.555 69.925 ;
        RECT 836.130 61.890 836.420 73.725 ;
        RECT 839.580 72.165 839.990 75.260 ;
        RECT 844.035 71.620 844.345 74.135 ;
        RECT 837.025 64.385 837.355 70.580 ;
        RECT 839.945 63.855 840.385 67.130 ;
        RECT 842.325 65.870 842.850 69.810 ;
        RECT 841.485 61.765 841.810 64.530 ;
        RECT 844.000 63.860 844.415 66.250 ;
        RECT 845.030 62.420 845.345 73.105 ;
        RECT 846.360 66.810 846.845 69.820 ;
        RECT 847.540 62.435 847.870 73.130 ;
        RECT 845.730 61.030 846.065 62.380 ;
        RECT 757.345 42.140 757.660 53.190 ;
        RECT 761.180 52.485 761.580 55.535 ;
        RECT 766.100 52.395 766.510 55.490 ;
        RECT 770.680 52.370 771.090 55.465 ;
        RECT 759.015 40.290 759.360 42.750 ;
        RECT 776.130 42.625 776.445 53.310 ;
        RECT 781.315 45.415 781.765 49.575 ;
        RECT 783.015 48.395 783.540 48.835 ;
        RECT 594.345 29.355 594.725 29.735 ;
        RECT 594.335 28.605 594.715 28.985 ;
        RECT 594.380 27.920 594.760 28.300 ;
        RECT 594.345 27.250 594.725 27.630 ;
        RECT 595.060 24.175 595.360 31.215 ;
        RECT 596.180 23.570 596.480 30.500 ;
        RECT 596.835 24.930 597.135 28.990 ;
        RECT 597.490 24.170 597.790 30.520 ;
        RECT 598.085 26.045 598.405 31.205 ;
        RECT 598.805 24.200 599.100 31.025 ;
        RECT 599.935 23.660 600.235 30.470 ;
        RECT 600.725 24.255 601.035 30.445 ;
        RECT 601.520 24.185 601.820 31.015 ;
        RECT 602.645 23.570 602.945 30.510 ;
        RECT 603.325 24.915 603.605 29.005 ;
        RECT 604.095 23.445 604.375 26.480 ;
        RECT 604.855 24.145 605.160 30.505 ;
        RECT 605.705 24.145 606.005 30.965 ;
        RECT 606.845 23.400 607.145 30.555 ;
        RECT 607.510 29.355 607.890 29.735 ;
        RECT 609.780 29.355 610.160 29.760 ;
        RECT 607.515 28.605 607.895 28.985 ;
        RECT 609.785 28.605 610.165 29.010 ;
        RECT 607.515 27.590 607.895 27.970 ;
        RECT 609.300 26.170 609.620 28.300 ;
        RECT 607.730 22.880 608.110 25.900 ;
        RECT 609.910 25.330 610.190 27.735 ;
        RECT 610.520 24.175 610.820 31.215 ;
        RECT 611.640 23.570 611.940 30.500 ;
        RECT 612.295 24.930 612.595 28.990 ;
        RECT 612.950 24.170 613.250 30.520 ;
        RECT 613.545 26.045 613.870 31.205 ;
        RECT 614.265 24.200 614.560 31.025 ;
        RECT 615.395 23.660 615.695 30.470 ;
        RECT 616.185 24.255 616.495 30.445 ;
        RECT 616.980 24.185 617.280 31.015 ;
        RECT 618.105 23.570 618.405 30.510 ;
        RECT 618.785 24.915 619.065 29.005 ;
        RECT 619.555 23.445 619.835 26.480 ;
        RECT 620.315 24.145 620.635 30.505 ;
        RECT 621.165 24.145 621.465 30.965 ;
        RECT 622.305 23.400 622.605 30.555 ;
        RECT 623.245 29.355 623.605 31.185 ;
        RECT 622.940 25.545 623.320 25.925 ;
        RECT 623.645 21.430 624.005 27.990 ;
        RECT 624.785 26.180 625.110 28.045 ;
        RECT 625.425 27.835 625.840 31.185 ;
        RECT 625.450 22.835 625.910 27.520 ;
        RECT 626.235 25.380 626.685 34.200 ;
        RECT 627.095 23.005 627.450 33.310 ;
        RECT 627.760 28.610 628.105 29.665 ;
        RECT 628.420 27.205 628.850 30.195 ;
        RECT 626.165 21.490 626.545 21.870 ;
        RECT 629.055 21.510 629.435 22.885 ;
        RECT 629.825 22.330 630.140 33.380 ;
        RECT 630.840 32.075 631.130 34.135 ;
        RECT 633.625 32.675 634.100 35.725 ;
        RECT 638.580 32.585 638.990 35.680 ;
        RECT 637.620 30.925 637.930 30.955 ;
        RECT 630.760 24.220 631.085 26.590 ;
        RECT 632.410 26.265 632.810 30.230 ;
        RECT 631.495 20.480 631.840 22.940 ;
        RECT 633.130 22.160 633.455 24.925 ;
        RECT 634.115 24.195 634.520 27.525 ;
        RECT 637.620 24.825 637.935 30.925 ;
        RECT 638.765 21.220 639.135 30.320 ;
        RECT 639.710 22.285 640.000 34.120 ;
        RECT 643.160 32.560 643.570 35.655 ;
        RECT 647.615 32.015 647.925 34.530 ;
        RECT 640.605 24.780 640.935 30.975 ;
        RECT 643.525 24.250 643.965 27.525 ;
        RECT 645.905 26.265 646.430 30.205 ;
        RECT 645.065 22.160 645.390 24.925 ;
        RECT 647.580 24.255 647.995 26.645 ;
        RECT 648.610 22.815 648.925 33.500 ;
        RECT 649.940 27.205 650.425 30.215 ;
        RECT 651.120 22.830 651.450 33.525 ;
        RECT 656.400 29.125 659.725 29.715 ;
        RECT 656.400 28.510 657.150 29.125 ;
        RECT 658.305 25.670 658.975 28.320 ;
        RECT 649.310 21.425 649.645 22.775 ;
        RECT 660.265 9.515 660.715 28.555 ;
        RECT 662.055 8.740 662.470 29.920 ;
        RECT 665.795 22.340 666.150 33.425 ;
        RECT 669.540 32.065 669.830 34.125 ;
        RECT 672.310 32.665 672.810 35.715 ;
        RECT 677.280 32.575 677.690 35.670 ;
        RECT 676.320 30.915 676.630 30.945 ;
        RECT 667.120 27.195 667.590 30.185 ;
        RECT 669.470 24.210 669.785 26.580 ;
        RECT 671.090 26.255 671.510 30.220 ;
        RECT 667.755 21.500 668.135 22.875 ;
        RECT 670.195 20.470 670.540 22.930 ;
        RECT 671.830 22.150 672.155 24.915 ;
        RECT 672.815 24.185 673.220 27.515 ;
        RECT 676.320 24.815 676.635 30.915 ;
        RECT 677.465 21.210 677.835 30.310 ;
        RECT 678.410 22.275 678.700 34.110 ;
        RECT 681.860 32.550 682.270 35.645 ;
        RECT 686.315 32.005 686.625 34.520 ;
        RECT 690.565 33.705 690.945 34.085 ;
        RECT 692.695 33.705 693.075 34.085 ;
        RECT 679.305 24.770 679.635 30.965 ;
        RECT 682.210 24.240 682.665 27.515 ;
        RECT 684.570 26.255 685.115 30.195 ;
        RECT 688.625 27.195 689.060 30.205 ;
        RECT 683.765 22.150 684.090 24.915 ;
        RECT 686.280 24.245 686.695 26.635 ;
        RECT 689.820 22.820 690.150 33.515 ;
        RECT 691.255 27.155 691.640 32.940 ;
        RECT 688.010 21.415 688.345 22.765 ;
        RECT 691.615 22.400 692.040 26.675 ;
        RECT 693.315 24.165 693.615 31.205 ;
        RECT 694.435 23.560 694.735 30.490 ;
        RECT 695.745 24.160 696.045 30.510 ;
        RECT 690.275 21.490 690.655 21.870 ;
        RECT 692.470 21.475 692.850 21.855 ;
        RECT 696.340 21.415 696.630 31.195 ;
        RECT 697.060 24.190 697.355 31.015 ;
        RECT 698.190 23.650 698.490 30.460 ;
        RECT 698.980 24.245 699.290 34.285 ;
        RECT 708.170 32.530 708.550 32.910 ;
        RECT 699.775 24.175 700.075 31.005 ;
        RECT 700.900 23.560 701.200 30.500 ;
        RECT 702.350 23.435 702.630 26.470 ;
        RECT 703.110 24.135 703.390 30.495 ;
        RECT 703.960 24.135 704.260 30.955 ;
        RECT 705.100 23.390 705.400 30.545 ;
        RECT 705.745 27.580 706.125 27.960 ;
        RECT 705.745 25.525 706.125 25.905 ;
        RECT 707.595 25.405 707.910 29.730 ;
        RECT 708.205 27.480 708.485 29.010 ;
        RECT 708.775 24.165 709.075 31.205 ;
        RECT 709.895 23.560 710.195 30.490 ;
        RECT 710.550 24.920 710.850 28.980 ;
        RECT 711.205 24.160 711.505 30.510 ;
        RECT 708.070 22.355 708.450 22.735 ;
        RECT 711.800 21.950 712.090 31.195 ;
        RECT 712.520 24.190 712.815 31.015 ;
        RECT 713.650 23.650 713.950 30.460 ;
        RECT 714.440 24.245 714.750 32.980 ;
        RECT 715.235 24.175 715.535 31.005 ;
        RECT 716.360 23.560 716.660 30.500 ;
        RECT 717.040 24.905 717.320 28.995 ;
        RECT 717.810 23.435 718.090 26.470 ;
        RECT 718.570 24.135 718.850 30.495 ;
        RECT 719.420 24.135 719.720 30.955 ;
        RECT 720.560 23.390 720.860 30.545 ;
        RECT 722.485 29.310 722.860 37.150 ;
        RECT 724.340 28.560 724.640 39.100 ;
        RECT 725.565 27.445 725.945 37.700 ;
        RECT 726.435 25.290 726.870 38.865 ;
        RECT 782.145 38.130 782.660 48.180 ;
        RECT 783.830 36.775 784.415 47.555 ;
        RECT 785.450 45.060 785.805 58.970 ;
        RECT 848.795 58.340 849.245 68.605 ;
        RECT 787.075 45.980 787.435 57.370 ;
        RECT 849.960 56.800 850.445 65.685 ;
        RECT 856.790 56.155 857.195 68.035 ;
        RECT 858.865 58.055 859.255 69.635 ;
        RECT 862.135 61.975 862.490 73.060 ;
        RECT 865.880 71.700 866.170 73.760 ;
        RECT 868.650 72.300 869.150 75.350 ;
        RECT 873.620 72.210 874.030 75.305 ;
        RECT 872.660 70.550 872.970 70.580 ;
        RECT 863.460 66.830 863.930 69.820 ;
        RECT 865.810 63.845 866.125 66.215 ;
        RECT 867.430 65.890 867.850 69.855 ;
        RECT 864.095 61.135 864.475 62.510 ;
        RECT 866.535 60.105 866.880 62.565 ;
        RECT 868.170 61.785 868.495 64.550 ;
        RECT 869.155 63.820 869.560 67.150 ;
        RECT 872.660 64.450 872.975 70.550 ;
        RECT 873.805 60.845 874.175 69.945 ;
        RECT 874.750 61.910 875.040 73.745 ;
        RECT 878.200 72.185 878.610 75.280 ;
        RECT 882.655 71.640 882.965 74.155 ;
        RECT 886.905 73.340 887.285 73.720 ;
        RECT 889.035 73.340 889.415 73.720 ;
        RECT 875.645 64.405 875.975 70.600 ;
        RECT 878.550 63.875 879.005 67.150 ;
        RECT 880.910 65.890 881.455 69.830 ;
        RECT 884.965 66.830 885.400 69.840 ;
        RECT 880.105 61.785 880.430 64.550 ;
        RECT 882.620 63.880 883.035 66.270 ;
        RECT 886.160 62.455 886.490 73.150 ;
        RECT 887.595 66.790 887.980 72.575 ;
        RECT 884.350 61.050 884.685 62.400 ;
        RECT 887.955 62.035 888.380 66.310 ;
        RECT 889.655 63.800 889.955 70.840 ;
        RECT 890.775 63.195 891.075 70.125 ;
        RECT 892.085 63.795 892.385 70.145 ;
        RECT 886.615 61.125 886.995 61.505 ;
        RECT 888.810 61.110 889.190 61.490 ;
        RECT 892.680 61.050 892.970 70.830 ;
        RECT 893.400 63.825 893.695 70.650 ;
        RECT 894.530 63.285 894.830 70.095 ;
        RECT 895.320 63.880 895.630 73.920 ;
        RECT 904.510 72.165 904.890 72.545 ;
        RECT 896.115 63.810 896.415 70.640 ;
        RECT 897.240 63.195 897.540 70.135 ;
        RECT 898.690 63.070 898.970 66.105 ;
        RECT 899.450 63.770 899.730 70.130 ;
        RECT 900.300 63.770 900.600 70.590 ;
        RECT 901.440 63.025 901.740 70.180 ;
        RECT 902.085 67.215 902.465 67.595 ;
        RECT 902.085 65.160 902.465 65.540 ;
        RECT 903.935 65.040 904.250 69.365 ;
        RECT 904.545 67.115 904.825 68.645 ;
        RECT 905.115 63.800 905.415 70.840 ;
        RECT 906.235 63.195 906.535 70.125 ;
        RECT 906.890 64.555 907.190 68.615 ;
        RECT 907.545 63.795 907.845 70.145 ;
        RECT 904.410 61.990 904.790 62.370 ;
        RECT 908.140 61.585 908.430 70.830 ;
        RECT 908.860 63.825 909.155 70.650 ;
        RECT 909.990 63.285 910.290 70.095 ;
        RECT 910.780 63.880 911.090 72.615 ;
        RECT 911.575 63.810 911.875 70.640 ;
        RECT 912.700 63.195 913.000 70.135 ;
        RECT 913.380 64.540 913.660 68.630 ;
        RECT 914.150 63.070 914.430 66.105 ;
        RECT 914.910 63.770 915.190 70.130 ;
        RECT 915.760 63.770 916.060 70.590 ;
        RECT 916.900 63.025 917.200 70.180 ;
        RECT 918.980 68.900 919.355 77.180 ;
        RECT 920.725 68.060 921.025 79.170 ;
        RECT 921.950 67.065 922.330 77.320 ;
        RECT 922.820 64.910 923.255 78.485 ;
        RECT 978.530 77.685 979.045 87.735 ;
        RECT 980.215 76.330 980.800 87.110 ;
        RECT 982.000 84.585 982.355 98.375 ;
        RECT 1045.345 97.745 1045.795 108.235 ;
        RECT 983.625 85.490 983.985 96.775 ;
        RECT 1046.510 96.205 1046.995 105.365 ;
        RECT 1052.970 96.015 1053.375 107.545 ;
        RECT 1055.045 97.915 1055.435 109.015 ;
        RECT 1058.450 101.445 1058.805 112.530 ;
        RECT 1062.195 111.170 1062.485 113.230 ;
        RECT 1064.965 111.770 1065.465 114.820 ;
        RECT 1069.935 111.680 1070.345 114.775 ;
        RECT 1068.975 110.020 1069.285 110.050 ;
        RECT 1059.775 106.300 1060.245 109.290 ;
        RECT 1062.125 103.315 1062.440 105.685 ;
        RECT 1063.745 105.360 1064.165 109.325 ;
        RECT 1060.410 100.605 1060.790 101.980 ;
        RECT 1062.850 99.575 1063.195 102.035 ;
        RECT 1064.485 101.255 1064.810 104.020 ;
        RECT 1065.470 103.290 1065.875 106.620 ;
        RECT 1068.975 103.920 1069.290 110.020 ;
        RECT 1070.120 100.315 1070.490 109.415 ;
        RECT 1071.065 101.380 1071.355 113.215 ;
        RECT 1074.515 111.655 1074.925 114.750 ;
        RECT 1078.970 111.110 1079.280 113.625 ;
        RECT 1083.220 112.810 1083.600 113.190 ;
        RECT 1085.350 112.810 1085.730 113.190 ;
        RECT 1071.960 103.875 1072.290 110.070 ;
        RECT 1074.865 103.345 1075.320 106.620 ;
        RECT 1077.225 105.360 1077.770 109.300 ;
        RECT 1081.280 106.300 1081.715 109.310 ;
        RECT 1076.420 101.255 1076.745 104.020 ;
        RECT 1078.935 103.350 1079.350 105.740 ;
        RECT 1082.475 101.925 1082.805 112.620 ;
        RECT 1083.910 106.260 1084.295 112.045 ;
        RECT 1080.665 100.520 1081.000 101.870 ;
        RECT 1084.270 101.505 1084.695 105.780 ;
        RECT 1085.970 103.270 1086.270 110.310 ;
        RECT 1087.090 102.665 1087.390 109.595 ;
        RECT 1088.400 103.265 1088.700 109.615 ;
        RECT 1082.930 100.595 1083.310 100.975 ;
        RECT 1085.125 100.580 1085.505 100.960 ;
        RECT 1088.995 100.520 1089.285 110.300 ;
        RECT 1089.715 103.295 1090.010 110.120 ;
        RECT 1090.845 102.755 1091.145 109.565 ;
        RECT 1091.635 103.350 1091.945 113.390 ;
        RECT 1100.825 111.635 1101.205 112.015 ;
        RECT 1092.430 103.280 1092.730 110.110 ;
        RECT 1093.555 102.665 1093.855 109.605 ;
        RECT 1095.005 102.540 1095.285 105.575 ;
        RECT 1095.765 103.240 1096.045 109.600 ;
        RECT 1096.615 103.240 1096.915 110.060 ;
        RECT 1097.755 102.495 1098.055 109.650 ;
        RECT 1098.400 106.685 1098.780 107.065 ;
        RECT 1098.400 104.630 1098.780 105.010 ;
        RECT 1100.250 104.510 1100.565 108.835 ;
        RECT 1100.860 106.585 1101.140 108.115 ;
        RECT 1101.430 103.270 1101.730 110.310 ;
        RECT 1102.550 102.665 1102.850 109.595 ;
        RECT 1103.205 104.025 1103.505 108.085 ;
        RECT 1103.860 103.265 1104.160 109.615 ;
        RECT 1100.725 101.460 1101.105 101.840 ;
        RECT 1104.455 101.055 1104.745 110.300 ;
        RECT 1105.175 103.295 1105.470 110.120 ;
        RECT 1106.305 102.755 1106.605 109.565 ;
        RECT 1107.095 103.350 1107.405 112.085 ;
        RECT 1107.890 103.280 1108.190 110.110 ;
        RECT 1109.015 102.665 1109.315 109.605 ;
        RECT 1109.695 104.010 1109.975 108.100 ;
        RECT 1110.465 102.540 1110.745 105.575 ;
        RECT 1111.225 103.240 1111.505 109.600 ;
        RECT 1112.075 103.240 1112.375 110.060 ;
        RECT 1113.215 102.495 1113.515 109.650 ;
        RECT 1115.420 108.420 1115.795 116.620 ;
        RECT 1117.165 107.615 1117.465 118.610 ;
        RECT 1118.275 106.535 1118.655 116.790 ;
        RECT 1119.145 104.380 1119.580 117.955 ;
        RECT 1175.000 117.235 1175.515 127.285 ;
        RECT 1176.685 115.880 1177.270 126.660 ;
        RECT 1178.175 124.150 1178.530 138.205 ;
        RECT 1241.520 137.575 1241.970 147.690 ;
        RECT 1179.800 124.955 1180.160 136.605 ;
        RECT 1242.685 136.035 1243.170 144.790 ;
        RECT 1249.290 135.410 1249.695 146.940 ;
        RECT 1251.365 137.310 1251.755 148.410 ;
        RECT 1254.635 140.885 1254.990 151.970 ;
        RECT 1255.960 145.740 1256.430 148.730 ;
        RECT 1256.595 140.045 1256.975 141.420 ;
        RECT 1257.365 140.865 1257.680 151.915 ;
        RECT 1258.380 150.610 1258.670 152.670 ;
        RECT 1261.150 151.210 1261.650 154.260 ;
        RECT 1266.120 151.120 1266.530 154.215 ;
        RECT 1265.160 149.460 1265.470 149.490 ;
        RECT 1258.310 142.755 1258.625 145.125 ;
        RECT 1259.930 144.800 1260.350 148.765 ;
        RECT 1259.035 139.015 1259.380 141.475 ;
        RECT 1260.670 140.695 1260.995 143.460 ;
        RECT 1261.655 142.730 1262.060 146.060 ;
        RECT 1265.160 143.360 1265.475 149.460 ;
        RECT 1266.305 139.755 1266.675 148.855 ;
        RECT 1267.250 140.820 1267.540 152.655 ;
        RECT 1270.700 151.095 1271.110 154.190 ;
        RECT 1275.155 150.550 1275.465 153.065 ;
        RECT 1279.405 152.250 1279.785 152.630 ;
        RECT 1281.535 152.250 1281.915 152.630 ;
        RECT 1268.145 143.315 1268.475 149.510 ;
        RECT 1271.050 142.785 1271.505 146.060 ;
        RECT 1273.410 144.800 1273.955 148.740 ;
        RECT 1272.605 140.695 1272.930 143.460 ;
        RECT 1275.120 142.790 1275.535 145.180 ;
        RECT 1276.150 141.350 1276.465 152.035 ;
        RECT 1277.465 145.740 1277.900 148.750 ;
        RECT 1278.660 141.365 1278.990 152.060 ;
        RECT 1279.340 147.110 1279.760 147.570 ;
        RECT 1280.095 145.700 1280.480 151.485 ;
        RECT 1280.840 147.105 1281.260 147.565 ;
        RECT 1279.475 144.220 1279.855 144.600 ;
        RECT 1276.850 139.960 1277.185 141.310 ;
        RECT 1280.455 140.945 1280.880 145.220 ;
        RECT 1281.540 144.195 1281.850 148.315 ;
        RECT 1282.155 142.710 1282.455 149.750 ;
        RECT 1283.275 142.105 1283.575 149.035 ;
        RECT 1283.930 143.465 1284.230 147.525 ;
        RECT 1284.585 142.705 1284.885 149.055 ;
        RECT 1279.115 140.035 1279.495 140.415 ;
        RECT 1281.310 140.020 1281.690 140.400 ;
        RECT 1285.180 139.960 1285.470 149.740 ;
        RECT 1285.900 142.735 1286.195 149.560 ;
        RECT 1287.030 142.195 1287.330 149.005 ;
        RECT 1287.820 142.790 1288.130 152.830 ;
        RECT 1288.615 142.720 1288.915 149.550 ;
        RECT 1289.740 142.105 1290.040 149.045 ;
        RECT 1290.420 143.450 1290.700 147.540 ;
        RECT 1291.190 141.980 1291.470 145.015 ;
        RECT 1291.950 142.680 1292.230 149.040 ;
        RECT 1292.800 142.680 1293.100 149.500 ;
        RECT 1293.940 141.935 1294.240 149.090 ;
        RECT 1294.610 147.890 1294.905 153.260 ;
        RECT 1295.185 147.060 1295.490 152.535 ;
        RECT 1297.010 151.075 1297.390 151.455 ;
        RECT 1294.585 146.125 1294.965 146.505 ;
        RECT 1294.585 144.070 1294.965 144.450 ;
        RECT 1296.435 143.950 1296.750 148.275 ;
        RECT 1297.045 146.025 1297.325 147.555 ;
        RECT 1297.615 142.710 1297.915 149.750 ;
        RECT 1299.390 143.465 1299.690 147.525 ;
        RECT 1296.910 140.900 1297.290 141.280 ;
        RECT 1300.640 140.495 1300.930 149.740 ;
        RECT 1302.490 142.195 1302.790 149.005 ;
        RECT 1303.280 142.790 1303.590 151.525 ;
        RECT 1304.075 142.720 1304.375 149.550 ;
        RECT 1305.880 143.450 1306.160 147.540 ;
        RECT 1306.650 141.980 1306.930 145.015 ;
        RECT 1309.400 141.935 1309.700 149.090 ;
        RECT 1311.440 147.830 1311.815 156.030 ;
        RECT 1313.185 147.025 1313.485 158.020 ;
        RECT 1183.640 128.270 1184.020 128.650 ;
        RECT 1183.630 127.520 1184.010 127.900 ;
        RECT 1183.675 126.835 1184.055 127.215 ;
        RECT 1183.640 126.165 1184.020 126.545 ;
        RECT 1184.355 123.090 1184.655 130.130 ;
        RECT 1185.475 122.485 1185.775 129.415 ;
        RECT 1186.130 123.845 1186.430 127.905 ;
        RECT 1186.785 123.085 1187.085 129.435 ;
        RECT 1187.380 124.960 1187.700 130.120 ;
        RECT 1188.100 123.115 1188.395 129.940 ;
        RECT 1189.230 122.575 1189.530 129.385 ;
        RECT 1190.020 123.170 1190.330 129.360 ;
        RECT 1190.815 123.100 1191.115 129.930 ;
        RECT 1191.940 122.485 1192.240 129.425 ;
        RECT 1192.620 123.830 1192.900 127.920 ;
        RECT 1193.390 122.360 1193.670 125.395 ;
        RECT 1194.150 123.060 1194.455 129.420 ;
        RECT 1195.000 123.060 1195.300 129.880 ;
        RECT 1196.140 122.315 1196.440 129.470 ;
        RECT 1196.805 128.270 1197.185 128.650 ;
        RECT 1199.075 128.270 1199.455 128.675 ;
        RECT 1196.810 127.520 1197.190 127.900 ;
        RECT 1199.080 127.520 1199.460 127.925 ;
        RECT 1196.810 126.505 1197.190 126.885 ;
        RECT 1198.595 125.085 1198.915 127.215 ;
        RECT 1197.025 121.795 1197.405 124.815 ;
        RECT 1199.205 124.245 1199.485 126.650 ;
        RECT 1199.815 123.090 1200.115 130.130 ;
        RECT 1200.935 122.485 1201.235 129.415 ;
        RECT 1201.590 123.845 1201.890 127.905 ;
        RECT 1202.245 123.085 1202.545 129.435 ;
        RECT 1202.840 124.960 1203.165 130.120 ;
        RECT 1203.560 123.115 1203.855 129.940 ;
        RECT 1204.690 122.575 1204.990 129.385 ;
        RECT 1205.480 123.170 1205.790 129.360 ;
        RECT 1206.275 123.100 1206.575 129.930 ;
        RECT 1207.400 122.485 1207.700 129.425 ;
        RECT 1208.080 123.830 1208.360 127.920 ;
        RECT 1208.850 122.360 1209.130 125.395 ;
        RECT 1209.610 123.060 1209.930 129.420 ;
        RECT 1210.460 123.060 1210.760 129.880 ;
        RECT 1211.600 122.315 1211.900 129.470 ;
        RECT 1212.540 128.270 1212.900 130.100 ;
        RECT 1212.235 124.460 1212.615 124.840 ;
        RECT 1212.940 120.345 1213.300 126.905 ;
        RECT 1214.080 125.095 1214.405 126.960 ;
        RECT 1214.720 126.750 1215.135 130.100 ;
        RECT 1214.745 121.750 1215.205 126.435 ;
        RECT 1215.530 124.295 1215.980 133.115 ;
        RECT 1216.390 121.920 1216.745 132.225 ;
        RECT 1217.055 127.525 1217.400 128.580 ;
        RECT 1217.715 126.120 1218.145 129.110 ;
        RECT 1215.460 120.405 1215.840 120.785 ;
        RECT 1218.350 120.425 1218.730 121.800 ;
        RECT 1219.120 121.245 1219.435 132.295 ;
        RECT 1220.135 130.990 1220.425 133.050 ;
        RECT 1222.920 131.590 1223.395 134.640 ;
        RECT 1227.875 131.500 1228.285 134.595 ;
        RECT 1226.915 129.840 1227.225 129.870 ;
        RECT 1220.055 123.135 1220.380 125.505 ;
        RECT 1221.705 125.180 1222.105 129.145 ;
        RECT 1220.790 119.395 1221.135 121.855 ;
        RECT 1222.425 121.075 1222.750 123.840 ;
        RECT 1223.410 123.110 1223.815 126.440 ;
        RECT 1226.915 123.740 1227.230 129.840 ;
        RECT 1228.060 120.135 1228.430 129.235 ;
        RECT 1229.005 121.200 1229.295 133.035 ;
        RECT 1232.455 131.475 1232.865 134.570 ;
        RECT 1236.910 130.930 1237.220 133.445 ;
        RECT 1229.900 123.695 1230.230 129.890 ;
        RECT 1232.820 123.165 1233.260 126.440 ;
        RECT 1235.200 125.180 1235.725 129.120 ;
        RECT 1234.360 121.075 1234.685 123.840 ;
        RECT 1236.875 123.170 1237.290 125.560 ;
        RECT 1237.905 121.730 1238.220 132.415 ;
        RECT 1239.235 126.120 1239.720 129.130 ;
        RECT 1240.415 121.745 1240.745 132.440 ;
        RECT 1238.605 120.340 1238.940 121.690 ;
        RECT 1150.025 101.405 1150.340 112.455 ;
        RECT 1153.860 111.750 1154.260 114.800 ;
        RECT 1158.780 111.660 1159.190 114.755 ;
        RECT 1163.360 111.635 1163.770 114.730 ;
        RECT 1151.695 99.555 1152.040 102.015 ;
        RECT 1168.810 101.890 1169.125 112.575 ;
        RECT 1173.995 104.680 1174.445 108.840 ;
        RECT 1175.695 107.660 1176.220 108.100 ;
        RECT 986.975 88.720 987.355 89.100 ;
        RECT 986.965 87.970 987.345 88.350 ;
        RECT 987.010 87.285 987.390 87.665 ;
        RECT 986.975 86.615 987.355 86.995 ;
        RECT 987.690 83.540 987.990 90.580 ;
        RECT 988.810 82.935 989.110 89.865 ;
        RECT 989.465 84.295 989.765 88.355 ;
        RECT 990.120 83.535 990.420 89.885 ;
        RECT 990.715 85.410 991.035 90.570 ;
        RECT 991.435 83.565 991.730 90.390 ;
        RECT 992.565 83.025 992.865 89.835 ;
        RECT 993.355 83.620 993.665 89.810 ;
        RECT 994.150 83.550 994.450 90.380 ;
        RECT 995.275 82.935 995.575 89.875 ;
        RECT 995.955 84.280 996.235 88.370 ;
        RECT 996.725 82.810 997.005 85.845 ;
        RECT 997.485 83.510 997.790 89.870 ;
        RECT 998.335 83.510 998.635 90.330 ;
        RECT 999.475 82.765 999.775 89.920 ;
        RECT 1000.140 88.720 1000.520 89.100 ;
        RECT 1002.410 88.720 1002.790 89.125 ;
        RECT 1000.145 87.970 1000.525 88.350 ;
        RECT 1002.415 87.970 1002.795 88.375 ;
        RECT 1000.145 86.955 1000.525 87.335 ;
        RECT 1001.930 85.535 1002.250 87.665 ;
        RECT 1000.360 82.245 1000.740 85.265 ;
        RECT 1002.540 84.695 1002.820 87.100 ;
        RECT 1003.150 83.540 1003.450 90.580 ;
        RECT 1004.270 82.935 1004.570 89.865 ;
        RECT 1004.925 84.295 1005.225 88.355 ;
        RECT 1005.580 83.535 1005.880 89.885 ;
        RECT 1006.175 85.410 1006.500 90.570 ;
        RECT 1006.895 83.565 1007.190 90.390 ;
        RECT 1008.025 83.025 1008.325 89.835 ;
        RECT 1008.815 83.620 1009.125 89.810 ;
        RECT 1009.610 83.550 1009.910 90.380 ;
        RECT 1010.735 82.935 1011.035 89.875 ;
        RECT 1011.415 84.280 1011.695 88.370 ;
        RECT 1012.185 82.810 1012.465 85.845 ;
        RECT 1012.945 83.510 1013.265 89.870 ;
        RECT 1013.795 83.510 1014.095 90.330 ;
        RECT 1014.935 82.765 1015.235 89.920 ;
        RECT 1015.875 88.720 1016.235 90.550 ;
        RECT 1015.570 84.910 1015.950 85.290 ;
        RECT 1016.275 80.795 1016.635 87.355 ;
        RECT 1017.415 85.545 1017.740 87.410 ;
        RECT 1018.055 87.200 1018.470 90.550 ;
        RECT 1018.080 82.200 1018.540 86.885 ;
        RECT 1018.865 84.745 1019.315 93.565 ;
        RECT 1019.725 82.370 1020.080 92.675 ;
        RECT 1020.390 87.975 1020.735 89.030 ;
        RECT 1021.050 86.570 1021.480 89.560 ;
        RECT 1018.795 80.855 1019.175 81.235 ;
        RECT 1021.685 80.875 1022.065 82.250 ;
        RECT 1022.455 81.695 1022.770 92.745 ;
        RECT 1023.470 91.440 1023.760 93.500 ;
        RECT 1026.255 92.040 1026.730 95.090 ;
        RECT 1031.210 91.950 1031.620 95.045 ;
        RECT 1030.250 90.290 1030.560 90.320 ;
        RECT 1023.390 83.585 1023.715 85.955 ;
        RECT 1025.040 85.630 1025.440 89.595 ;
        RECT 1024.125 79.845 1024.470 82.305 ;
        RECT 1025.760 81.525 1026.085 84.290 ;
        RECT 1026.745 83.560 1027.150 86.890 ;
        RECT 1030.250 84.190 1030.565 90.290 ;
        RECT 1031.395 80.585 1031.765 89.685 ;
        RECT 1032.340 81.650 1032.630 93.485 ;
        RECT 1035.790 91.925 1036.200 95.020 ;
        RECT 1040.245 91.380 1040.555 93.895 ;
        RECT 1033.235 84.145 1033.565 90.340 ;
        RECT 1036.155 83.615 1036.595 86.890 ;
        RECT 1038.535 85.630 1039.060 89.570 ;
        RECT 1037.695 81.525 1038.020 84.290 ;
        RECT 1040.210 83.620 1040.625 86.010 ;
        RECT 1041.240 82.180 1041.555 92.865 ;
        RECT 1042.570 86.570 1043.055 89.580 ;
        RECT 1043.750 82.195 1044.080 92.890 ;
        RECT 1041.940 80.790 1042.275 82.140 ;
        RECT 953.660 61.845 953.975 72.895 ;
        RECT 957.495 72.190 957.895 75.240 ;
        RECT 962.415 72.100 962.825 75.195 ;
        RECT 966.995 72.075 967.405 75.170 ;
        RECT 955.330 59.995 955.675 62.455 ;
        RECT 972.445 62.330 972.760 73.015 ;
        RECT 977.630 65.120 978.080 69.280 ;
        RECT 979.330 68.100 979.855 68.540 ;
        RECT 790.715 49.150 791.095 49.530 ;
        RECT 790.705 48.400 791.085 48.780 ;
        RECT 790.750 47.715 791.130 48.095 ;
        RECT 790.715 47.045 791.095 47.425 ;
        RECT 791.430 43.970 791.730 51.010 ;
        RECT 792.550 43.365 792.850 50.295 ;
        RECT 793.205 44.725 793.505 48.785 ;
        RECT 793.860 43.965 794.160 50.315 ;
        RECT 794.455 45.840 794.775 51.000 ;
        RECT 795.175 43.995 795.470 50.820 ;
        RECT 796.305 43.455 796.605 50.265 ;
        RECT 797.095 44.050 797.405 50.240 ;
        RECT 797.890 43.980 798.190 50.810 ;
        RECT 799.015 43.365 799.315 50.305 ;
        RECT 799.695 44.710 799.975 48.800 ;
        RECT 800.465 43.240 800.745 46.275 ;
        RECT 801.225 43.940 801.530 50.300 ;
        RECT 802.075 43.940 802.375 50.760 ;
        RECT 803.215 43.195 803.515 50.350 ;
        RECT 803.880 49.150 804.260 49.530 ;
        RECT 806.150 49.150 806.530 49.555 ;
        RECT 803.885 48.400 804.265 48.780 ;
        RECT 806.155 48.400 806.535 48.805 ;
        RECT 803.885 47.385 804.265 47.765 ;
        RECT 805.670 45.965 805.990 48.095 ;
        RECT 804.100 42.675 804.480 45.695 ;
        RECT 806.280 45.125 806.560 47.530 ;
        RECT 806.890 43.970 807.190 51.010 ;
        RECT 808.010 43.365 808.310 50.295 ;
        RECT 808.665 44.725 808.965 48.785 ;
        RECT 809.320 43.965 809.620 50.315 ;
        RECT 809.915 45.840 810.240 51.000 ;
        RECT 810.635 43.995 810.930 50.820 ;
        RECT 811.765 43.455 812.065 50.265 ;
        RECT 812.555 44.050 812.865 50.240 ;
        RECT 813.350 43.980 813.650 50.810 ;
        RECT 814.475 43.365 814.775 50.305 ;
        RECT 815.155 44.710 815.435 48.800 ;
        RECT 815.925 43.240 816.205 46.275 ;
        RECT 816.685 43.940 817.005 50.300 ;
        RECT 817.535 43.940 817.835 50.760 ;
        RECT 818.675 43.195 818.975 50.350 ;
        RECT 819.615 49.150 819.975 50.980 ;
        RECT 819.310 45.340 819.690 45.720 ;
        RECT 820.015 41.225 820.375 47.785 ;
        RECT 821.155 45.975 821.480 47.840 ;
        RECT 821.795 47.630 822.210 50.980 ;
        RECT 821.820 42.630 822.280 47.315 ;
        RECT 822.605 45.175 823.055 53.995 ;
        RECT 823.465 42.800 823.820 53.105 ;
        RECT 824.130 48.405 824.475 49.460 ;
        RECT 824.790 47.000 825.220 49.990 ;
        RECT 822.535 41.285 822.915 41.665 ;
        RECT 825.425 41.305 825.805 42.680 ;
        RECT 826.195 42.125 826.510 53.175 ;
        RECT 827.210 51.870 827.500 53.930 ;
        RECT 829.995 52.470 830.470 55.520 ;
        RECT 834.950 52.380 835.360 55.475 ;
        RECT 833.990 50.720 834.300 50.750 ;
        RECT 827.130 44.015 827.455 46.385 ;
        RECT 828.780 46.060 829.180 50.025 ;
        RECT 827.865 40.275 828.210 42.735 ;
        RECT 829.500 41.955 829.825 44.720 ;
        RECT 830.485 43.990 830.890 47.320 ;
        RECT 833.990 44.620 834.305 50.720 ;
        RECT 835.135 41.015 835.505 50.115 ;
        RECT 836.080 42.080 836.370 53.915 ;
        RECT 839.530 52.355 839.940 55.450 ;
        RECT 843.985 51.810 844.295 54.325 ;
        RECT 836.975 44.575 837.305 50.770 ;
        RECT 839.895 44.045 840.335 47.320 ;
        RECT 842.275 46.060 842.800 50.000 ;
        RECT 841.435 41.955 841.760 44.720 ;
        RECT 843.950 44.050 844.365 46.440 ;
        RECT 844.980 42.610 845.295 53.295 ;
        RECT 846.310 47.000 846.795 50.010 ;
        RECT 847.490 42.625 847.820 53.320 ;
        RECT 845.680 41.220 846.015 42.570 ;
        RECT 757.320 22.410 757.635 33.460 ;
        RECT 761.155 32.755 761.555 35.805 ;
        RECT 766.075 32.665 766.485 35.760 ;
        RECT 770.655 32.640 771.065 35.735 ;
        RECT 758.990 20.560 759.335 23.020 ;
        RECT 776.105 22.895 776.420 33.580 ;
        RECT 781.340 25.610 781.790 29.770 ;
        RECT 783.040 28.590 783.565 29.030 ;
        RECT 665.815 3.825 666.115 10.755 ;
        RECT 666.470 5.185 666.770 9.245 ;
        RECT 667.125 4.425 667.425 10.775 ;
        RECT 668.440 4.455 668.735 11.280 ;
        RECT 672.280 3.825 672.580 10.765 ;
        RECT 672.960 5.170 673.240 9.260 ;
        RECT 674.490 4.400 674.795 10.760 ;
        RECT 675.340 4.400 675.640 11.220 ;
        RECT 677.070 7.840 677.450 8.220 ;
        RECT 677.080 5.795 677.460 6.175 ;
        RECT 782.140 5.450 782.655 27.705 ;
        RECT 783.825 7.665 784.410 28.385 ;
        RECT 785.450 25.220 785.805 39.160 ;
        RECT 848.795 38.530 849.245 48.795 ;
        RECT 787.075 26.010 787.435 37.560 ;
        RECT 849.960 36.990 850.445 45.875 ;
        RECT 856.900 36.265 857.305 48.310 ;
        RECT 858.975 38.165 859.365 49.590 ;
        RECT 862.135 42.005 862.490 53.090 ;
        RECT 865.880 51.730 866.170 53.790 ;
        RECT 868.650 52.330 869.150 55.380 ;
        RECT 873.620 52.240 874.030 55.335 ;
        RECT 872.660 50.580 872.970 50.610 ;
        RECT 863.460 46.860 863.930 49.850 ;
        RECT 865.810 43.875 866.125 46.245 ;
        RECT 867.430 45.920 867.850 49.885 ;
        RECT 864.095 41.165 864.475 42.540 ;
        RECT 866.535 40.135 866.880 42.595 ;
        RECT 868.170 41.815 868.495 44.580 ;
        RECT 869.155 43.850 869.560 47.180 ;
        RECT 872.660 44.480 872.975 50.580 ;
        RECT 873.805 40.875 874.175 49.975 ;
        RECT 874.750 41.940 875.040 53.775 ;
        RECT 878.200 52.215 878.610 55.310 ;
        RECT 882.655 51.670 882.965 54.185 ;
        RECT 886.905 53.370 887.285 53.750 ;
        RECT 889.035 53.370 889.415 53.750 ;
        RECT 875.645 44.435 875.975 50.630 ;
        RECT 878.550 43.905 879.005 47.180 ;
        RECT 880.910 45.920 881.455 49.860 ;
        RECT 884.965 46.860 885.400 49.870 ;
        RECT 880.105 41.815 880.430 44.580 ;
        RECT 882.620 43.910 883.035 46.300 ;
        RECT 886.160 42.485 886.490 53.180 ;
        RECT 887.595 46.820 887.980 52.605 ;
        RECT 884.350 41.080 884.685 42.430 ;
        RECT 887.955 42.065 888.380 46.340 ;
        RECT 889.655 43.830 889.955 50.870 ;
        RECT 890.775 43.225 891.075 50.155 ;
        RECT 892.085 43.825 892.385 50.175 ;
        RECT 886.615 41.155 886.995 41.535 ;
        RECT 888.810 41.140 889.190 41.520 ;
        RECT 892.680 41.080 892.970 50.860 ;
        RECT 893.400 43.855 893.695 50.680 ;
        RECT 894.530 43.315 894.830 50.125 ;
        RECT 895.320 43.910 895.630 53.950 ;
        RECT 904.510 52.195 904.890 52.575 ;
        RECT 896.115 43.840 896.415 50.670 ;
        RECT 897.240 43.225 897.540 50.165 ;
        RECT 898.690 43.100 898.970 46.135 ;
        RECT 899.450 43.800 899.730 50.160 ;
        RECT 900.300 43.800 900.600 50.620 ;
        RECT 901.440 43.055 901.740 50.210 ;
        RECT 902.085 47.245 902.465 47.625 ;
        RECT 902.085 45.190 902.465 45.570 ;
        RECT 903.935 45.070 904.250 49.395 ;
        RECT 904.545 47.145 904.825 48.675 ;
        RECT 905.115 43.830 905.415 50.870 ;
        RECT 906.235 43.225 906.535 50.155 ;
        RECT 906.890 44.585 907.190 48.645 ;
        RECT 907.545 43.825 907.845 50.175 ;
        RECT 904.410 42.020 904.790 42.400 ;
        RECT 908.140 41.615 908.430 50.860 ;
        RECT 908.860 43.855 909.155 50.680 ;
        RECT 909.990 43.315 910.290 50.125 ;
        RECT 910.780 43.910 911.090 52.645 ;
        RECT 911.575 43.840 911.875 50.670 ;
        RECT 912.700 43.225 913.000 50.165 ;
        RECT 913.380 44.570 913.660 48.660 ;
        RECT 914.150 43.100 914.430 46.135 ;
        RECT 914.910 43.800 915.190 50.160 ;
        RECT 915.760 43.800 916.060 50.620 ;
        RECT 916.900 43.055 917.200 50.210 ;
        RECT 919.240 48.825 919.615 57.025 ;
        RECT 920.985 48.020 921.285 59.015 ;
        RECT 921.950 47.090 922.330 57.345 ;
        RECT 922.820 44.935 923.255 58.510 ;
        RECT 978.530 57.670 979.045 67.970 ;
        RECT 980.215 56.565 980.800 67.345 ;
        RECT 981.695 64.825 982.050 78.745 ;
        RECT 1045.040 78.115 1045.490 88.380 ;
        RECT 983.320 65.730 983.680 77.145 ;
        RECT 1046.205 76.575 1046.690 85.460 ;
        RECT 1052.870 76.310 1053.275 87.840 ;
        RECT 1054.945 78.210 1055.335 89.310 ;
        RECT 1058.370 81.690 1058.725 92.775 ;
        RECT 1062.115 91.415 1062.405 93.475 ;
        RECT 1064.885 92.015 1065.385 95.065 ;
        RECT 1069.855 91.925 1070.265 95.020 ;
        RECT 1068.895 90.265 1069.205 90.295 ;
        RECT 1059.695 86.545 1060.165 89.535 ;
        RECT 1062.045 83.560 1062.360 85.930 ;
        RECT 1063.665 85.605 1064.085 89.570 ;
        RECT 1060.330 80.850 1060.710 82.225 ;
        RECT 1062.770 79.820 1063.115 82.280 ;
        RECT 1064.405 81.500 1064.730 84.265 ;
        RECT 1065.390 83.535 1065.795 86.865 ;
        RECT 1068.895 84.165 1069.210 90.265 ;
        RECT 1070.040 80.560 1070.410 89.660 ;
        RECT 1070.985 81.625 1071.275 93.460 ;
        RECT 1074.435 91.900 1074.845 94.995 ;
        RECT 1078.890 91.355 1079.200 93.870 ;
        RECT 1083.140 93.055 1083.520 93.435 ;
        RECT 1085.270 93.055 1085.650 93.435 ;
        RECT 1071.880 84.120 1072.210 90.315 ;
        RECT 1074.785 83.590 1075.240 86.865 ;
        RECT 1077.145 85.605 1077.690 89.545 ;
        RECT 1081.200 86.545 1081.635 89.555 ;
        RECT 1076.340 81.500 1076.665 84.265 ;
        RECT 1078.855 83.595 1079.270 85.985 ;
        RECT 1082.395 82.170 1082.725 92.865 ;
        RECT 1083.830 86.505 1084.215 92.290 ;
        RECT 1080.585 80.765 1080.920 82.115 ;
        RECT 1084.190 81.750 1084.615 86.025 ;
        RECT 1085.890 83.515 1086.190 90.555 ;
        RECT 1087.010 82.910 1087.310 89.840 ;
        RECT 1088.320 83.510 1088.620 89.860 ;
        RECT 1082.850 80.840 1083.230 81.220 ;
        RECT 1085.045 80.825 1085.425 81.205 ;
        RECT 1088.915 80.765 1089.205 90.545 ;
        RECT 1089.635 83.540 1089.930 90.365 ;
        RECT 1090.765 83.000 1091.065 89.810 ;
        RECT 1091.555 83.595 1091.865 93.635 ;
        RECT 1100.745 91.880 1101.125 92.260 ;
        RECT 1092.350 83.525 1092.650 90.355 ;
        RECT 1093.475 82.910 1093.775 89.850 ;
        RECT 1094.925 82.785 1095.205 85.820 ;
        RECT 1095.685 83.485 1095.965 89.845 ;
        RECT 1096.535 83.485 1096.835 90.305 ;
        RECT 1097.675 82.740 1097.975 89.895 ;
        RECT 1098.320 86.930 1098.700 87.310 ;
        RECT 1098.320 84.875 1098.700 85.255 ;
        RECT 1100.170 84.755 1100.485 89.080 ;
        RECT 1100.780 86.830 1101.060 88.360 ;
        RECT 1101.350 83.515 1101.650 90.555 ;
        RECT 1102.470 82.910 1102.770 89.840 ;
        RECT 1103.125 84.270 1103.425 88.330 ;
        RECT 1103.780 83.510 1104.080 89.860 ;
        RECT 1100.645 81.705 1101.025 82.085 ;
        RECT 1104.375 81.300 1104.665 90.545 ;
        RECT 1105.095 83.540 1105.390 90.365 ;
        RECT 1106.225 83.000 1106.525 89.810 ;
        RECT 1107.015 83.595 1107.325 92.330 ;
        RECT 1107.810 83.525 1108.110 90.355 ;
        RECT 1108.935 82.910 1109.235 89.850 ;
        RECT 1109.615 84.255 1109.895 88.345 ;
        RECT 1110.385 82.785 1110.665 85.820 ;
        RECT 1111.145 83.485 1111.425 89.845 ;
        RECT 1111.995 83.485 1112.295 90.305 ;
        RECT 1113.135 82.740 1113.435 89.895 ;
        RECT 1115.420 88.600 1115.795 96.885 ;
        RECT 1117.165 87.880 1117.465 98.875 ;
        RECT 1118.275 86.780 1118.655 97.035 ;
        RECT 1119.145 84.625 1119.580 98.200 ;
        RECT 1174.850 97.400 1175.365 107.450 ;
        RECT 1176.535 96.045 1177.120 106.825 ;
        RECT 1178.385 104.375 1178.740 118.165 ;
        RECT 1241.730 117.535 1242.180 128.035 ;
        RECT 1180.010 105.230 1180.370 116.565 ;
        RECT 1242.895 115.995 1243.380 125.235 ;
        RECT 1249.310 115.750 1249.715 127.280 ;
        RECT 1251.385 117.650 1251.775 128.750 ;
        RECT 1254.790 121.240 1255.145 132.325 ;
        RECT 1256.115 126.095 1256.585 129.085 ;
        RECT 1256.750 120.400 1257.130 121.775 ;
        RECT 1257.520 121.220 1257.835 132.270 ;
        RECT 1258.535 130.965 1258.825 133.025 ;
        RECT 1261.305 131.565 1261.805 134.615 ;
        RECT 1266.275 131.475 1266.685 134.570 ;
        RECT 1265.315 129.815 1265.625 129.845 ;
        RECT 1258.465 123.110 1258.780 125.480 ;
        RECT 1260.085 125.155 1260.505 129.120 ;
        RECT 1259.190 119.370 1259.535 121.830 ;
        RECT 1260.825 121.050 1261.150 123.815 ;
        RECT 1261.810 123.085 1262.215 126.415 ;
        RECT 1265.315 123.715 1265.630 129.815 ;
        RECT 1266.460 120.110 1266.830 129.210 ;
        RECT 1267.405 121.175 1267.695 133.010 ;
        RECT 1270.855 131.450 1271.265 134.545 ;
        RECT 1275.310 130.905 1275.620 133.420 ;
        RECT 1279.560 132.605 1279.940 132.985 ;
        RECT 1281.690 132.605 1282.070 132.985 ;
        RECT 1268.300 123.670 1268.630 129.865 ;
        RECT 1271.205 123.140 1271.660 126.415 ;
        RECT 1273.565 125.155 1274.110 129.095 ;
        RECT 1272.760 121.050 1273.085 123.815 ;
        RECT 1275.275 123.145 1275.690 125.535 ;
        RECT 1276.305 121.705 1276.620 132.390 ;
        RECT 1277.620 126.095 1278.055 129.105 ;
        RECT 1278.815 121.720 1279.145 132.415 ;
        RECT 1279.495 127.465 1279.915 127.925 ;
        RECT 1280.250 126.055 1280.635 131.840 ;
        RECT 1280.995 127.460 1281.415 127.920 ;
        RECT 1279.630 124.575 1280.010 124.955 ;
        RECT 1277.005 120.315 1277.340 121.665 ;
        RECT 1280.610 121.300 1281.035 125.575 ;
        RECT 1281.695 124.550 1282.005 128.670 ;
        RECT 1282.310 123.065 1282.610 130.105 ;
        RECT 1283.430 122.460 1283.730 129.390 ;
        RECT 1284.085 123.820 1284.385 127.880 ;
        RECT 1284.740 123.060 1285.040 129.410 ;
        RECT 1279.270 120.390 1279.650 120.770 ;
        RECT 1281.465 120.375 1281.845 120.755 ;
        RECT 1285.335 120.315 1285.625 130.095 ;
        RECT 1286.055 123.090 1286.350 129.915 ;
        RECT 1287.185 122.550 1287.485 129.360 ;
        RECT 1287.975 123.145 1288.285 133.185 ;
        RECT 1288.770 123.075 1289.070 129.905 ;
        RECT 1289.895 122.460 1290.195 129.400 ;
        RECT 1290.575 123.805 1290.855 127.895 ;
        RECT 1291.345 122.335 1291.625 125.370 ;
        RECT 1292.105 123.035 1292.385 129.395 ;
        RECT 1292.955 123.035 1293.255 129.855 ;
        RECT 1294.095 122.290 1294.395 129.445 ;
        RECT 1294.765 128.245 1295.060 133.615 ;
        RECT 1295.340 127.415 1295.645 132.890 ;
        RECT 1297.165 131.430 1297.545 131.810 ;
        RECT 1294.740 126.480 1295.120 126.860 ;
        RECT 1294.740 124.425 1295.120 124.805 ;
        RECT 1296.590 124.305 1296.905 128.630 ;
        RECT 1297.200 126.380 1297.480 127.910 ;
        RECT 1297.770 123.065 1298.070 130.105 ;
        RECT 1299.545 123.820 1299.845 127.880 ;
        RECT 1297.065 121.255 1297.445 121.635 ;
        RECT 1300.795 120.850 1301.085 130.095 ;
        RECT 1302.645 122.550 1302.945 129.360 ;
        RECT 1303.435 123.145 1303.745 131.880 ;
        RECT 1304.230 123.075 1304.530 129.905 ;
        RECT 1306.035 123.805 1306.315 127.895 ;
        RECT 1306.805 122.335 1307.085 125.370 ;
        RECT 1309.555 122.290 1309.855 129.445 ;
        RECT 1311.740 128.080 1312.115 136.280 ;
        RECT 1313.485 127.275 1313.785 138.270 ;
        RECT 1183.445 108.430 1183.825 108.810 ;
        RECT 1183.435 107.680 1183.815 108.060 ;
        RECT 1183.480 106.995 1183.860 107.375 ;
        RECT 1183.445 106.325 1183.825 106.705 ;
        RECT 1184.160 103.250 1184.460 110.290 ;
        RECT 1185.280 102.645 1185.580 109.575 ;
        RECT 1185.935 104.005 1186.235 108.065 ;
        RECT 1186.590 103.245 1186.890 109.595 ;
        RECT 1187.185 105.120 1187.505 110.280 ;
        RECT 1187.905 103.275 1188.200 110.100 ;
        RECT 1189.035 102.735 1189.335 109.545 ;
        RECT 1189.825 103.330 1190.135 109.520 ;
        RECT 1190.620 103.260 1190.920 110.090 ;
        RECT 1191.745 102.645 1192.045 109.585 ;
        RECT 1192.425 103.990 1192.705 108.080 ;
        RECT 1193.195 102.520 1193.475 105.555 ;
        RECT 1193.955 103.220 1194.260 109.580 ;
        RECT 1194.805 103.220 1195.105 110.040 ;
        RECT 1195.945 102.475 1196.245 109.630 ;
        RECT 1196.610 108.430 1196.990 108.810 ;
        RECT 1198.880 108.430 1199.260 108.835 ;
        RECT 1196.615 107.680 1196.995 108.060 ;
        RECT 1198.885 107.680 1199.265 108.085 ;
        RECT 1196.615 106.665 1196.995 107.045 ;
        RECT 1198.400 105.245 1198.720 107.375 ;
        RECT 1196.830 101.955 1197.210 104.975 ;
        RECT 1199.010 104.405 1199.290 106.810 ;
        RECT 1199.620 103.250 1199.920 110.290 ;
        RECT 1200.740 102.645 1201.040 109.575 ;
        RECT 1201.395 104.005 1201.695 108.065 ;
        RECT 1202.050 103.245 1202.350 109.595 ;
        RECT 1202.645 105.120 1202.970 110.280 ;
        RECT 1203.365 103.275 1203.660 110.100 ;
        RECT 1204.495 102.735 1204.795 109.545 ;
        RECT 1205.285 103.330 1205.595 109.520 ;
        RECT 1206.080 103.260 1206.380 110.090 ;
        RECT 1207.205 102.645 1207.505 109.585 ;
        RECT 1207.885 103.990 1208.165 108.080 ;
        RECT 1208.655 102.520 1208.935 105.555 ;
        RECT 1209.415 103.220 1209.735 109.580 ;
        RECT 1210.265 103.220 1210.565 110.040 ;
        RECT 1211.405 102.475 1211.705 109.630 ;
        RECT 1212.345 108.430 1212.705 110.260 ;
        RECT 1212.040 104.620 1212.420 105.000 ;
        RECT 1212.745 100.505 1213.105 107.065 ;
        RECT 1213.885 105.255 1214.210 107.120 ;
        RECT 1214.525 106.910 1214.940 110.260 ;
        RECT 1214.550 101.910 1215.010 106.595 ;
        RECT 1215.335 104.455 1215.785 113.275 ;
        RECT 1216.195 102.080 1216.550 112.385 ;
        RECT 1216.860 107.685 1217.205 108.740 ;
        RECT 1217.520 106.280 1217.950 109.270 ;
        RECT 1215.265 100.565 1215.645 100.945 ;
        RECT 1218.155 100.585 1218.535 101.960 ;
        RECT 1218.925 101.405 1219.240 112.455 ;
        RECT 1219.940 111.150 1220.230 113.210 ;
        RECT 1222.725 111.750 1223.200 114.800 ;
        RECT 1227.680 111.660 1228.090 114.755 ;
        RECT 1226.720 110.000 1227.030 110.030 ;
        RECT 1219.860 103.295 1220.185 105.665 ;
        RECT 1221.510 105.340 1221.910 109.305 ;
        RECT 1220.595 99.555 1220.940 102.015 ;
        RECT 1222.230 101.235 1222.555 104.000 ;
        RECT 1223.215 103.270 1223.620 106.600 ;
        RECT 1226.720 103.900 1227.035 110.000 ;
        RECT 1227.865 100.295 1228.235 109.395 ;
        RECT 1228.810 101.360 1229.100 113.195 ;
        RECT 1232.260 111.635 1232.670 114.730 ;
        RECT 1236.715 111.090 1237.025 113.605 ;
        RECT 1229.705 103.855 1230.035 110.050 ;
        RECT 1232.625 103.325 1233.065 106.600 ;
        RECT 1235.005 105.340 1235.530 109.280 ;
        RECT 1234.165 101.235 1234.490 104.000 ;
        RECT 1236.680 103.330 1237.095 105.720 ;
        RECT 1237.710 101.890 1238.025 112.575 ;
        RECT 1239.040 106.280 1239.525 109.290 ;
        RECT 1240.220 101.905 1240.550 112.600 ;
        RECT 1238.410 100.500 1238.745 101.850 ;
        RECT 1150.055 81.680 1150.370 92.730 ;
        RECT 1153.890 92.025 1154.290 95.075 ;
        RECT 1158.810 91.935 1159.220 95.030 ;
        RECT 1163.390 91.910 1163.800 95.005 ;
        RECT 1151.725 79.830 1152.070 82.290 ;
        RECT 1168.840 82.165 1169.155 92.850 ;
        RECT 1174.025 84.955 1174.475 89.115 ;
        RECT 1175.725 87.935 1176.250 88.375 ;
        RECT 987.105 68.960 987.485 69.340 ;
        RECT 987.095 68.210 987.475 68.590 ;
        RECT 987.140 67.525 987.520 67.905 ;
        RECT 987.105 66.855 987.485 67.235 ;
        RECT 987.820 63.780 988.120 70.820 ;
        RECT 988.940 63.175 989.240 70.105 ;
        RECT 989.595 64.535 989.895 68.595 ;
        RECT 990.250 63.775 990.550 70.125 ;
        RECT 990.845 65.650 991.165 70.810 ;
        RECT 991.565 63.805 991.860 70.630 ;
        RECT 992.695 63.265 992.995 70.075 ;
        RECT 993.485 63.860 993.795 70.050 ;
        RECT 994.280 63.790 994.580 70.620 ;
        RECT 995.405 63.175 995.705 70.115 ;
        RECT 996.085 64.520 996.365 68.610 ;
        RECT 996.855 63.050 997.135 66.085 ;
        RECT 997.615 63.750 997.920 70.110 ;
        RECT 998.465 63.750 998.765 70.570 ;
        RECT 999.605 63.005 999.905 70.160 ;
        RECT 1000.270 68.960 1000.650 69.340 ;
        RECT 1002.540 68.960 1002.920 69.365 ;
        RECT 1000.275 68.210 1000.655 68.590 ;
        RECT 1002.545 68.210 1002.925 68.615 ;
        RECT 1000.275 67.195 1000.655 67.575 ;
        RECT 1002.060 65.775 1002.380 67.905 ;
        RECT 1000.490 62.485 1000.870 65.505 ;
        RECT 1002.670 64.935 1002.950 67.340 ;
        RECT 1003.280 63.780 1003.580 70.820 ;
        RECT 1004.400 63.175 1004.700 70.105 ;
        RECT 1005.055 64.535 1005.355 68.595 ;
        RECT 1005.710 63.775 1006.010 70.125 ;
        RECT 1006.305 65.650 1006.630 70.810 ;
        RECT 1007.025 63.805 1007.320 70.630 ;
        RECT 1008.155 63.265 1008.455 70.075 ;
        RECT 1008.945 63.860 1009.255 70.050 ;
        RECT 1009.740 63.790 1010.040 70.620 ;
        RECT 1010.865 63.175 1011.165 70.115 ;
        RECT 1011.545 64.520 1011.825 68.610 ;
        RECT 1012.315 63.050 1012.595 66.085 ;
        RECT 1013.075 63.750 1013.395 70.110 ;
        RECT 1013.925 63.750 1014.225 70.570 ;
        RECT 1015.065 63.005 1015.365 70.160 ;
        RECT 1016.005 68.960 1016.365 70.790 ;
        RECT 1015.700 65.150 1016.080 65.530 ;
        RECT 1016.405 61.035 1016.765 67.595 ;
        RECT 1017.545 65.785 1017.870 67.650 ;
        RECT 1018.185 67.440 1018.600 70.790 ;
        RECT 1018.210 62.440 1018.670 67.125 ;
        RECT 1018.995 64.985 1019.445 73.805 ;
        RECT 1019.855 62.610 1020.210 72.915 ;
        RECT 1020.520 68.215 1020.865 69.270 ;
        RECT 1021.180 66.810 1021.610 69.800 ;
        RECT 1018.925 61.095 1019.305 61.475 ;
        RECT 1021.815 61.115 1022.195 62.490 ;
        RECT 1022.585 61.935 1022.900 72.985 ;
        RECT 1023.600 71.680 1023.890 73.740 ;
        RECT 1026.385 72.280 1026.860 75.330 ;
        RECT 1031.340 72.190 1031.750 75.285 ;
        RECT 1030.380 70.530 1030.690 70.560 ;
        RECT 1023.520 63.825 1023.845 66.195 ;
        RECT 1025.170 65.870 1025.570 69.835 ;
        RECT 1024.255 60.085 1024.600 62.545 ;
        RECT 1025.890 61.765 1026.215 64.530 ;
        RECT 1026.875 63.800 1027.280 67.130 ;
        RECT 1030.380 64.430 1030.695 70.530 ;
        RECT 1031.525 60.825 1031.895 69.925 ;
        RECT 1032.470 61.890 1032.760 73.725 ;
        RECT 1035.920 72.165 1036.330 75.260 ;
        RECT 1040.375 71.620 1040.685 74.135 ;
        RECT 1033.365 64.385 1033.695 70.580 ;
        RECT 1036.285 63.855 1036.725 67.130 ;
        RECT 1038.665 65.870 1039.190 69.810 ;
        RECT 1037.825 61.765 1038.150 64.530 ;
        RECT 1040.340 63.860 1040.755 66.250 ;
        RECT 1041.370 62.420 1041.685 73.105 ;
        RECT 1042.700 66.810 1043.185 69.820 ;
        RECT 1043.880 62.435 1044.210 73.130 ;
        RECT 1042.070 61.030 1042.405 62.380 ;
        RECT 953.730 42.125 954.045 53.175 ;
        RECT 957.565 52.470 957.965 55.520 ;
        RECT 962.485 52.380 962.895 55.475 ;
        RECT 967.065 52.355 967.475 55.450 ;
        RECT 955.400 40.275 955.745 42.735 ;
        RECT 972.515 42.610 972.830 53.295 ;
        RECT 977.700 45.400 978.150 49.560 ;
        RECT 979.400 48.380 979.925 48.820 ;
        RECT 790.685 29.355 791.065 29.735 ;
        RECT 790.675 28.605 791.055 28.985 ;
        RECT 790.720 27.920 791.100 28.300 ;
        RECT 790.685 27.250 791.065 27.630 ;
        RECT 791.400 24.175 791.700 31.215 ;
        RECT 792.520 23.570 792.820 30.500 ;
        RECT 793.175 24.930 793.475 28.990 ;
        RECT 793.830 24.170 794.130 30.520 ;
        RECT 794.425 26.045 794.745 31.205 ;
        RECT 795.145 24.200 795.440 31.025 ;
        RECT 796.275 23.660 796.575 30.470 ;
        RECT 797.065 24.255 797.375 30.445 ;
        RECT 797.860 24.185 798.160 31.015 ;
        RECT 798.985 23.570 799.285 30.510 ;
        RECT 799.665 24.915 799.945 29.005 ;
        RECT 800.435 23.445 800.715 26.480 ;
        RECT 801.195 24.145 801.500 30.505 ;
        RECT 802.045 24.145 802.345 30.965 ;
        RECT 803.185 23.400 803.485 30.555 ;
        RECT 803.850 29.355 804.230 29.735 ;
        RECT 806.120 29.355 806.500 29.760 ;
        RECT 803.855 28.605 804.235 28.985 ;
        RECT 806.125 28.605 806.505 29.010 ;
        RECT 803.855 27.590 804.235 27.970 ;
        RECT 805.640 26.170 805.960 28.300 ;
        RECT 804.070 22.880 804.450 25.900 ;
        RECT 806.250 25.330 806.530 27.735 ;
        RECT 806.860 24.175 807.160 31.215 ;
        RECT 807.980 23.570 808.280 30.500 ;
        RECT 808.635 24.930 808.935 28.990 ;
        RECT 809.290 24.170 809.590 30.520 ;
        RECT 809.885 26.045 810.210 31.205 ;
        RECT 810.605 24.200 810.900 31.025 ;
        RECT 811.735 23.660 812.035 30.470 ;
        RECT 812.525 24.255 812.835 30.445 ;
        RECT 813.320 24.185 813.620 31.015 ;
        RECT 814.445 23.570 814.745 30.510 ;
        RECT 815.125 24.915 815.405 29.005 ;
        RECT 815.895 23.445 816.175 26.480 ;
        RECT 816.655 24.145 816.975 30.505 ;
        RECT 817.505 24.145 817.805 30.965 ;
        RECT 818.645 23.400 818.945 30.555 ;
        RECT 819.585 29.355 819.945 31.185 ;
        RECT 819.280 25.545 819.660 25.925 ;
        RECT 819.985 21.430 820.345 27.990 ;
        RECT 821.125 26.180 821.450 28.045 ;
        RECT 821.765 27.835 822.180 31.185 ;
        RECT 821.790 22.835 822.250 27.520 ;
        RECT 822.575 25.380 823.025 34.200 ;
        RECT 823.435 23.005 823.790 33.310 ;
        RECT 824.100 28.610 824.445 29.665 ;
        RECT 824.760 27.205 825.190 30.195 ;
        RECT 822.505 21.490 822.885 21.870 ;
        RECT 825.395 21.510 825.775 22.885 ;
        RECT 826.165 22.330 826.480 33.380 ;
        RECT 827.180 32.075 827.470 34.135 ;
        RECT 829.965 32.675 830.440 35.725 ;
        RECT 834.920 32.585 835.330 35.680 ;
        RECT 833.960 30.925 834.270 30.955 ;
        RECT 827.100 24.220 827.425 26.590 ;
        RECT 828.750 26.265 829.150 30.230 ;
        RECT 827.835 20.480 828.180 22.940 ;
        RECT 829.470 22.160 829.795 24.925 ;
        RECT 830.455 24.195 830.860 27.525 ;
        RECT 833.960 24.825 834.275 30.925 ;
        RECT 835.105 21.220 835.475 30.320 ;
        RECT 836.050 22.285 836.340 34.120 ;
        RECT 839.500 32.560 839.910 35.655 ;
        RECT 843.955 32.015 844.265 34.530 ;
        RECT 836.945 24.780 837.275 30.975 ;
        RECT 839.865 24.250 840.305 27.525 ;
        RECT 842.245 26.265 842.770 30.205 ;
        RECT 841.405 22.160 841.730 24.925 ;
        RECT 843.920 24.255 844.335 26.645 ;
        RECT 844.950 22.815 845.265 33.500 ;
        RECT 846.280 27.205 846.765 30.215 ;
        RECT 847.460 22.830 847.790 33.525 ;
        RECT 852.740 29.125 856.065 29.715 ;
        RECT 852.740 28.510 853.490 29.125 ;
        RECT 854.645 25.670 855.315 28.320 ;
        RECT 845.650 21.425 845.985 22.775 ;
        RECT 856.605 9.515 857.055 28.555 ;
        RECT 858.395 8.740 858.810 29.920 ;
        RECT 862.135 22.340 862.490 33.425 ;
        RECT 865.880 32.065 866.170 34.125 ;
        RECT 868.650 32.665 869.150 35.715 ;
        RECT 873.620 32.575 874.030 35.670 ;
        RECT 872.660 30.915 872.970 30.945 ;
        RECT 863.460 27.195 863.930 30.185 ;
        RECT 865.810 24.210 866.125 26.580 ;
        RECT 867.430 26.255 867.850 30.220 ;
        RECT 864.095 21.500 864.475 22.875 ;
        RECT 866.535 20.470 866.880 22.930 ;
        RECT 868.170 22.150 868.495 24.915 ;
        RECT 869.155 24.185 869.560 27.515 ;
        RECT 872.660 24.815 872.975 30.915 ;
        RECT 873.805 21.210 874.175 30.310 ;
        RECT 874.750 22.275 875.040 34.110 ;
        RECT 878.200 32.550 878.610 35.645 ;
        RECT 882.655 32.005 882.965 34.520 ;
        RECT 886.905 33.705 887.285 34.085 ;
        RECT 889.035 33.705 889.415 34.085 ;
        RECT 875.645 24.770 875.975 30.965 ;
        RECT 878.550 24.240 879.005 27.515 ;
        RECT 880.910 26.255 881.455 30.195 ;
        RECT 884.965 27.195 885.400 30.205 ;
        RECT 880.105 22.150 880.430 24.915 ;
        RECT 882.620 24.245 883.035 26.635 ;
        RECT 886.160 22.820 886.490 33.515 ;
        RECT 887.595 27.155 887.980 32.940 ;
        RECT 884.350 21.415 884.685 22.765 ;
        RECT 887.955 22.400 888.380 26.675 ;
        RECT 889.655 24.165 889.955 31.205 ;
        RECT 890.775 23.560 891.075 30.490 ;
        RECT 892.085 24.160 892.385 30.510 ;
        RECT 886.615 21.490 886.995 21.870 ;
        RECT 888.810 21.475 889.190 21.855 ;
        RECT 892.680 21.415 892.970 31.195 ;
        RECT 893.400 24.190 893.695 31.015 ;
        RECT 894.530 23.650 894.830 30.460 ;
        RECT 895.320 24.245 895.630 34.285 ;
        RECT 904.510 32.530 904.890 32.910 ;
        RECT 896.115 24.175 896.415 31.005 ;
        RECT 897.240 23.560 897.540 30.500 ;
        RECT 898.690 23.435 898.970 26.470 ;
        RECT 899.450 24.135 899.730 30.495 ;
        RECT 900.300 24.135 900.600 30.955 ;
        RECT 901.440 23.390 901.740 30.545 ;
        RECT 902.085 27.580 902.465 27.960 ;
        RECT 902.085 25.525 902.465 25.905 ;
        RECT 903.935 25.405 904.250 29.730 ;
        RECT 904.545 27.480 904.825 29.010 ;
        RECT 905.115 24.165 905.415 31.205 ;
        RECT 906.235 23.560 906.535 30.490 ;
        RECT 906.890 24.920 907.190 28.980 ;
        RECT 907.545 24.160 907.845 30.510 ;
        RECT 904.410 22.355 904.790 22.735 ;
        RECT 908.140 21.950 908.430 31.195 ;
        RECT 908.860 24.190 909.155 31.015 ;
        RECT 909.990 23.650 910.290 30.460 ;
        RECT 910.780 24.245 911.090 32.980 ;
        RECT 911.575 24.175 911.875 31.005 ;
        RECT 912.700 23.560 913.000 30.500 ;
        RECT 913.380 24.905 913.660 28.995 ;
        RECT 914.150 23.435 914.430 26.470 ;
        RECT 914.910 24.135 915.190 30.495 ;
        RECT 915.760 24.135 916.060 30.955 ;
        RECT 916.900 23.390 917.200 30.545 ;
        RECT 918.825 29.310 919.200 37.150 ;
        RECT 920.680 28.560 920.980 39.100 ;
        RECT 921.950 27.430 922.330 37.685 ;
        RECT 922.820 25.275 923.255 38.850 ;
        RECT 978.530 38.115 979.045 48.165 ;
        RECT 980.215 36.760 980.800 47.540 ;
        RECT 981.790 45.060 982.145 58.970 ;
        RECT 1045.135 58.340 1045.585 68.605 ;
        RECT 983.415 45.980 983.775 57.370 ;
        RECT 1046.300 56.800 1046.785 65.685 ;
        RECT 1053.130 56.155 1053.535 68.035 ;
        RECT 1055.205 58.055 1055.595 69.635 ;
        RECT 1058.475 61.975 1058.830 73.060 ;
        RECT 1062.220 71.700 1062.510 73.760 ;
        RECT 1064.990 72.300 1065.490 75.350 ;
        RECT 1069.960 72.210 1070.370 75.305 ;
        RECT 1069.000 70.550 1069.310 70.580 ;
        RECT 1059.800 66.830 1060.270 69.820 ;
        RECT 1062.150 63.845 1062.465 66.215 ;
        RECT 1063.770 65.890 1064.190 69.855 ;
        RECT 1060.435 61.135 1060.815 62.510 ;
        RECT 1062.875 60.105 1063.220 62.565 ;
        RECT 1064.510 61.785 1064.835 64.550 ;
        RECT 1065.495 63.820 1065.900 67.150 ;
        RECT 1069.000 64.450 1069.315 70.550 ;
        RECT 1070.145 60.845 1070.515 69.945 ;
        RECT 1071.090 61.910 1071.380 73.745 ;
        RECT 1074.540 72.185 1074.950 75.280 ;
        RECT 1078.995 71.640 1079.305 74.155 ;
        RECT 1083.245 73.340 1083.625 73.720 ;
        RECT 1085.375 73.340 1085.755 73.720 ;
        RECT 1071.985 64.405 1072.315 70.600 ;
        RECT 1074.890 63.875 1075.345 67.150 ;
        RECT 1077.250 65.890 1077.795 69.830 ;
        RECT 1081.305 66.830 1081.740 69.840 ;
        RECT 1076.445 61.785 1076.770 64.550 ;
        RECT 1078.960 63.880 1079.375 66.270 ;
        RECT 1082.500 62.455 1082.830 73.150 ;
        RECT 1083.935 66.790 1084.320 72.575 ;
        RECT 1080.690 61.050 1081.025 62.400 ;
        RECT 1084.295 62.035 1084.720 66.310 ;
        RECT 1085.995 63.800 1086.295 70.840 ;
        RECT 1087.115 63.195 1087.415 70.125 ;
        RECT 1088.425 63.795 1088.725 70.145 ;
        RECT 1082.955 61.125 1083.335 61.505 ;
        RECT 1085.150 61.110 1085.530 61.490 ;
        RECT 1089.020 61.050 1089.310 70.830 ;
        RECT 1089.740 63.825 1090.035 70.650 ;
        RECT 1090.870 63.285 1091.170 70.095 ;
        RECT 1091.660 63.880 1091.970 73.920 ;
        RECT 1100.850 72.165 1101.230 72.545 ;
        RECT 1092.455 63.810 1092.755 70.640 ;
        RECT 1093.580 63.195 1093.880 70.135 ;
        RECT 1095.030 63.070 1095.310 66.105 ;
        RECT 1095.790 63.770 1096.070 70.130 ;
        RECT 1096.640 63.770 1096.940 70.590 ;
        RECT 1097.780 63.025 1098.080 70.180 ;
        RECT 1098.425 67.215 1098.805 67.595 ;
        RECT 1098.425 65.160 1098.805 65.540 ;
        RECT 1100.275 65.040 1100.590 69.365 ;
        RECT 1100.885 67.115 1101.165 68.645 ;
        RECT 1101.455 63.800 1101.755 70.840 ;
        RECT 1102.575 63.195 1102.875 70.125 ;
        RECT 1103.230 64.555 1103.530 68.615 ;
        RECT 1103.885 63.795 1104.185 70.145 ;
        RECT 1100.750 61.990 1101.130 62.370 ;
        RECT 1104.480 61.585 1104.770 70.830 ;
        RECT 1105.200 63.825 1105.495 70.650 ;
        RECT 1106.330 63.285 1106.630 70.095 ;
        RECT 1107.120 63.880 1107.430 72.615 ;
        RECT 1107.915 63.810 1108.215 70.640 ;
        RECT 1109.040 63.195 1109.340 70.135 ;
        RECT 1109.720 64.540 1110.000 68.630 ;
        RECT 1110.490 63.070 1110.770 66.105 ;
        RECT 1111.250 63.770 1111.530 70.130 ;
        RECT 1112.100 63.770 1112.400 70.590 ;
        RECT 1113.240 63.025 1113.540 70.180 ;
        RECT 1115.320 68.900 1115.695 77.180 ;
        RECT 1117.065 68.060 1117.365 79.170 ;
        RECT 1118.275 67.070 1118.655 77.325 ;
        RECT 1119.145 64.915 1119.580 78.490 ;
        RECT 1174.855 77.690 1175.370 87.740 ;
        RECT 1176.540 76.335 1177.125 87.115 ;
        RECT 1178.340 84.585 1178.695 98.375 ;
        RECT 1241.685 97.745 1242.135 108.235 ;
        RECT 1179.965 85.490 1180.325 96.775 ;
        RECT 1242.850 96.205 1243.335 105.365 ;
        RECT 1249.310 96.015 1249.715 107.545 ;
        RECT 1251.385 97.915 1251.775 109.015 ;
        RECT 1254.790 101.445 1255.145 112.530 ;
        RECT 1256.115 106.300 1256.585 109.290 ;
        RECT 1256.750 100.605 1257.130 101.980 ;
        RECT 1257.520 101.425 1257.835 112.475 ;
        RECT 1258.535 111.170 1258.825 113.230 ;
        RECT 1261.305 111.770 1261.805 114.820 ;
        RECT 1266.275 111.680 1266.685 114.775 ;
        RECT 1265.315 110.020 1265.625 110.050 ;
        RECT 1258.465 103.315 1258.780 105.685 ;
        RECT 1260.085 105.360 1260.505 109.325 ;
        RECT 1259.190 99.575 1259.535 102.035 ;
        RECT 1260.825 101.255 1261.150 104.020 ;
        RECT 1261.810 103.290 1262.215 106.620 ;
        RECT 1265.315 103.920 1265.630 110.020 ;
        RECT 1266.460 100.315 1266.830 109.415 ;
        RECT 1267.405 101.380 1267.695 113.215 ;
        RECT 1270.855 111.655 1271.265 114.750 ;
        RECT 1275.310 111.110 1275.620 113.625 ;
        RECT 1279.560 112.810 1279.940 113.190 ;
        RECT 1281.690 112.810 1282.070 113.190 ;
        RECT 1268.300 103.875 1268.630 110.070 ;
        RECT 1271.205 103.345 1271.660 106.620 ;
        RECT 1273.565 105.360 1274.110 109.300 ;
        RECT 1272.760 101.255 1273.085 104.020 ;
        RECT 1275.275 103.350 1275.690 105.740 ;
        RECT 1276.305 101.910 1276.620 112.595 ;
        RECT 1277.620 106.300 1278.055 109.310 ;
        RECT 1278.815 101.925 1279.145 112.620 ;
        RECT 1279.495 107.670 1279.915 108.130 ;
        RECT 1280.250 106.260 1280.635 112.045 ;
        RECT 1280.995 107.665 1281.415 108.125 ;
        RECT 1279.630 104.780 1280.010 105.160 ;
        RECT 1277.005 100.520 1277.340 101.870 ;
        RECT 1280.610 101.505 1281.035 105.780 ;
        RECT 1281.695 104.755 1282.005 108.875 ;
        RECT 1282.310 103.270 1282.610 110.310 ;
        RECT 1283.430 102.665 1283.730 109.595 ;
        RECT 1284.085 104.025 1284.385 108.085 ;
        RECT 1284.740 103.265 1285.040 109.615 ;
        RECT 1279.270 100.595 1279.650 100.975 ;
        RECT 1281.465 100.580 1281.845 100.960 ;
        RECT 1285.335 100.520 1285.625 110.300 ;
        RECT 1286.055 103.295 1286.350 110.120 ;
        RECT 1287.185 102.755 1287.485 109.565 ;
        RECT 1287.975 103.350 1288.285 113.390 ;
        RECT 1288.770 103.280 1289.070 110.110 ;
        RECT 1289.895 102.665 1290.195 109.605 ;
        RECT 1290.575 104.010 1290.855 108.100 ;
        RECT 1291.345 102.540 1291.625 105.575 ;
        RECT 1292.105 103.240 1292.385 109.600 ;
        RECT 1292.955 103.240 1293.255 110.060 ;
        RECT 1294.095 102.495 1294.395 109.650 ;
        RECT 1294.765 108.450 1295.060 113.820 ;
        RECT 1295.340 107.620 1295.645 113.095 ;
        RECT 1297.165 111.635 1297.545 112.015 ;
        RECT 1294.740 106.685 1295.120 107.065 ;
        RECT 1294.740 104.630 1295.120 105.010 ;
        RECT 1296.590 104.510 1296.905 108.835 ;
        RECT 1297.200 106.585 1297.480 108.115 ;
        RECT 1297.770 103.270 1298.070 110.310 ;
        RECT 1299.545 104.025 1299.845 108.085 ;
        RECT 1297.065 101.460 1297.445 101.840 ;
        RECT 1300.795 101.055 1301.085 110.300 ;
        RECT 1302.645 102.755 1302.945 109.565 ;
        RECT 1303.435 103.350 1303.745 112.085 ;
        RECT 1304.230 103.280 1304.530 110.110 ;
        RECT 1306.035 104.010 1306.315 108.100 ;
        RECT 1306.805 102.540 1307.085 105.575 ;
        RECT 1309.555 102.495 1309.855 109.650 ;
        RECT 1311.760 108.420 1312.135 116.620 ;
        RECT 1313.505 107.615 1313.805 118.610 ;
        RECT 1183.315 88.720 1183.695 89.100 ;
        RECT 1183.305 87.970 1183.685 88.350 ;
        RECT 1183.350 87.285 1183.730 87.665 ;
        RECT 1183.315 86.615 1183.695 86.995 ;
        RECT 1184.030 83.540 1184.330 90.580 ;
        RECT 1185.150 82.935 1185.450 89.865 ;
        RECT 1185.805 84.295 1186.105 88.355 ;
        RECT 1186.460 83.535 1186.760 89.885 ;
        RECT 1187.055 85.410 1187.375 90.570 ;
        RECT 1187.775 83.565 1188.070 90.390 ;
        RECT 1188.905 83.025 1189.205 89.835 ;
        RECT 1189.695 83.620 1190.005 89.810 ;
        RECT 1190.490 83.550 1190.790 90.380 ;
        RECT 1191.615 82.935 1191.915 89.875 ;
        RECT 1192.295 84.280 1192.575 88.370 ;
        RECT 1193.065 82.810 1193.345 85.845 ;
        RECT 1193.825 83.510 1194.130 89.870 ;
        RECT 1194.675 83.510 1194.975 90.330 ;
        RECT 1195.815 82.765 1196.115 89.920 ;
        RECT 1196.480 88.720 1196.860 89.100 ;
        RECT 1198.750 88.720 1199.130 89.125 ;
        RECT 1196.485 87.970 1196.865 88.350 ;
        RECT 1198.755 87.970 1199.135 88.375 ;
        RECT 1196.485 86.955 1196.865 87.335 ;
        RECT 1198.270 85.535 1198.590 87.665 ;
        RECT 1196.700 82.245 1197.080 85.265 ;
        RECT 1198.880 84.695 1199.160 87.100 ;
        RECT 1199.490 83.540 1199.790 90.580 ;
        RECT 1200.610 82.935 1200.910 89.865 ;
        RECT 1201.265 84.295 1201.565 88.355 ;
        RECT 1201.920 83.535 1202.220 89.885 ;
        RECT 1202.515 85.410 1202.840 90.570 ;
        RECT 1203.235 83.565 1203.530 90.390 ;
        RECT 1204.365 83.025 1204.665 89.835 ;
        RECT 1205.155 83.620 1205.465 89.810 ;
        RECT 1205.950 83.550 1206.250 90.380 ;
        RECT 1207.075 82.935 1207.375 89.875 ;
        RECT 1207.755 84.280 1208.035 88.370 ;
        RECT 1208.525 82.810 1208.805 85.845 ;
        RECT 1209.285 83.510 1209.605 89.870 ;
        RECT 1210.135 83.510 1210.435 90.330 ;
        RECT 1211.275 82.765 1211.575 89.920 ;
        RECT 1212.215 88.720 1212.575 90.550 ;
        RECT 1211.910 84.910 1212.290 85.290 ;
        RECT 1212.615 80.795 1212.975 87.355 ;
        RECT 1213.755 85.545 1214.080 87.410 ;
        RECT 1214.395 87.200 1214.810 90.550 ;
        RECT 1214.420 82.200 1214.880 86.885 ;
        RECT 1215.205 84.745 1215.655 93.565 ;
        RECT 1216.065 82.370 1216.420 92.675 ;
        RECT 1216.730 87.975 1217.075 89.030 ;
        RECT 1217.390 86.570 1217.820 89.560 ;
        RECT 1215.135 80.855 1215.515 81.235 ;
        RECT 1218.025 80.875 1218.405 82.250 ;
        RECT 1218.795 81.695 1219.110 92.745 ;
        RECT 1219.810 91.440 1220.100 93.500 ;
        RECT 1222.595 92.040 1223.070 95.090 ;
        RECT 1227.550 91.950 1227.960 95.045 ;
        RECT 1226.590 90.290 1226.900 90.320 ;
        RECT 1219.730 83.585 1220.055 85.955 ;
        RECT 1221.380 85.630 1221.780 89.595 ;
        RECT 1220.465 79.845 1220.810 82.305 ;
        RECT 1222.100 81.525 1222.425 84.290 ;
        RECT 1223.085 83.560 1223.490 86.890 ;
        RECT 1226.590 84.190 1226.905 90.290 ;
        RECT 1227.735 80.585 1228.105 89.685 ;
        RECT 1228.680 81.650 1228.970 93.485 ;
        RECT 1232.130 91.925 1232.540 95.020 ;
        RECT 1236.585 91.380 1236.895 93.895 ;
        RECT 1229.575 84.145 1229.905 90.340 ;
        RECT 1232.495 83.615 1232.935 86.890 ;
        RECT 1234.875 85.630 1235.400 89.570 ;
        RECT 1234.035 81.525 1234.360 84.290 ;
        RECT 1236.550 83.620 1236.965 86.010 ;
        RECT 1237.580 82.180 1237.895 92.865 ;
        RECT 1238.910 86.570 1239.395 89.580 ;
        RECT 1240.090 82.195 1240.420 92.890 ;
        RECT 1238.280 80.790 1238.615 82.140 ;
        RECT 1149.985 61.850 1150.300 72.900 ;
        RECT 1153.820 72.195 1154.220 75.245 ;
        RECT 1158.740 72.105 1159.150 75.200 ;
        RECT 1163.320 72.080 1163.730 75.175 ;
        RECT 1151.655 60.000 1152.000 62.460 ;
        RECT 1168.770 62.335 1169.085 73.020 ;
        RECT 1173.955 65.125 1174.405 69.285 ;
        RECT 1175.655 68.105 1176.180 68.545 ;
        RECT 987.055 49.150 987.435 49.530 ;
        RECT 987.045 48.400 987.425 48.780 ;
        RECT 987.090 47.715 987.470 48.095 ;
        RECT 987.055 47.045 987.435 47.425 ;
        RECT 987.770 43.970 988.070 51.010 ;
        RECT 988.890 43.365 989.190 50.295 ;
        RECT 989.545 44.725 989.845 48.785 ;
        RECT 990.200 43.965 990.500 50.315 ;
        RECT 990.795 45.840 991.115 51.000 ;
        RECT 991.515 43.995 991.810 50.820 ;
        RECT 992.645 43.455 992.945 50.265 ;
        RECT 993.435 44.050 993.745 50.240 ;
        RECT 994.230 43.980 994.530 50.810 ;
        RECT 995.355 43.365 995.655 50.305 ;
        RECT 996.035 44.710 996.315 48.800 ;
        RECT 996.805 43.240 997.085 46.275 ;
        RECT 997.565 43.940 997.870 50.300 ;
        RECT 998.415 43.940 998.715 50.760 ;
        RECT 999.555 43.195 999.855 50.350 ;
        RECT 1000.220 49.150 1000.600 49.530 ;
        RECT 1002.490 49.150 1002.870 49.555 ;
        RECT 1000.225 48.400 1000.605 48.780 ;
        RECT 1002.495 48.400 1002.875 48.805 ;
        RECT 1000.225 47.385 1000.605 47.765 ;
        RECT 1002.010 45.965 1002.330 48.095 ;
        RECT 1000.440 42.675 1000.820 45.695 ;
        RECT 1002.620 45.125 1002.900 47.530 ;
        RECT 1003.230 43.970 1003.530 51.010 ;
        RECT 1004.350 43.365 1004.650 50.295 ;
        RECT 1005.005 44.725 1005.305 48.785 ;
        RECT 1005.660 43.965 1005.960 50.315 ;
        RECT 1006.255 45.840 1006.580 51.000 ;
        RECT 1006.975 43.995 1007.270 50.820 ;
        RECT 1008.105 43.455 1008.405 50.265 ;
        RECT 1008.895 44.050 1009.205 50.240 ;
        RECT 1009.690 43.980 1009.990 50.810 ;
        RECT 1010.815 43.365 1011.115 50.305 ;
        RECT 1011.495 44.710 1011.775 48.800 ;
        RECT 1012.265 43.240 1012.545 46.275 ;
        RECT 1013.025 43.940 1013.345 50.300 ;
        RECT 1013.875 43.940 1014.175 50.760 ;
        RECT 1015.015 43.195 1015.315 50.350 ;
        RECT 1015.955 49.150 1016.315 50.980 ;
        RECT 1015.650 45.340 1016.030 45.720 ;
        RECT 1016.355 41.225 1016.715 47.785 ;
        RECT 1017.495 45.975 1017.820 47.840 ;
        RECT 1018.135 47.630 1018.550 50.980 ;
        RECT 1018.160 42.630 1018.620 47.315 ;
        RECT 1018.945 45.175 1019.395 53.995 ;
        RECT 1019.805 42.800 1020.160 53.105 ;
        RECT 1020.470 48.405 1020.815 49.460 ;
        RECT 1021.130 47.000 1021.560 49.990 ;
        RECT 1018.875 41.285 1019.255 41.665 ;
        RECT 1021.765 41.305 1022.145 42.680 ;
        RECT 1022.535 42.125 1022.850 53.175 ;
        RECT 1023.550 51.870 1023.840 53.930 ;
        RECT 1026.335 52.470 1026.810 55.520 ;
        RECT 1031.290 52.380 1031.700 55.475 ;
        RECT 1030.330 50.720 1030.640 50.750 ;
        RECT 1023.470 44.015 1023.795 46.385 ;
        RECT 1025.120 46.060 1025.520 50.025 ;
        RECT 1024.205 40.275 1024.550 42.735 ;
        RECT 1025.840 41.955 1026.165 44.720 ;
        RECT 1026.825 43.990 1027.230 47.320 ;
        RECT 1030.330 44.620 1030.645 50.720 ;
        RECT 1031.475 41.015 1031.845 50.115 ;
        RECT 1032.420 42.080 1032.710 53.915 ;
        RECT 1035.870 52.355 1036.280 55.450 ;
        RECT 1040.325 51.810 1040.635 54.325 ;
        RECT 1033.315 44.575 1033.645 50.770 ;
        RECT 1036.235 44.045 1036.675 47.320 ;
        RECT 1038.615 46.060 1039.140 50.000 ;
        RECT 1037.775 41.955 1038.100 44.720 ;
        RECT 1040.290 44.050 1040.705 46.440 ;
        RECT 1041.320 42.610 1041.635 53.295 ;
        RECT 1042.650 47.000 1043.135 50.010 ;
        RECT 1043.830 42.625 1044.160 53.320 ;
        RECT 1042.020 41.220 1042.355 42.570 ;
        RECT 953.705 22.395 954.020 33.445 ;
        RECT 957.540 32.740 957.940 35.790 ;
        RECT 962.460 32.650 962.870 35.745 ;
        RECT 967.040 32.625 967.450 35.720 ;
        RECT 955.375 20.545 955.720 23.005 ;
        RECT 972.490 22.880 972.805 33.565 ;
        RECT 977.725 25.595 978.175 29.755 ;
        RECT 979.425 28.575 979.950 29.015 ;
        RECT 862.155 3.825 862.455 10.755 ;
        RECT 862.810 5.185 863.110 9.245 ;
        RECT 863.465 4.425 863.765 10.775 ;
        RECT 864.780 4.455 865.075 11.280 ;
        RECT 868.620 3.825 868.920 10.765 ;
        RECT 869.300 5.170 869.580 9.260 ;
        RECT 870.830 4.400 871.135 10.760 ;
        RECT 871.680 4.400 871.980 11.220 ;
        RECT 873.410 7.840 873.790 8.220 ;
        RECT 873.420 5.795 873.800 6.175 ;
        RECT 978.525 5.435 979.040 27.755 ;
        RECT 980.210 7.650 980.795 28.410 ;
        RECT 981.790 25.220 982.145 39.160 ;
        RECT 1045.135 38.530 1045.585 48.795 ;
        RECT 983.415 26.010 983.775 37.560 ;
        RECT 1046.300 36.990 1046.785 45.875 ;
        RECT 1053.240 36.265 1053.645 48.310 ;
        RECT 1055.315 38.165 1055.705 49.590 ;
        RECT 1058.475 42.005 1058.830 53.090 ;
        RECT 1062.220 51.730 1062.510 53.790 ;
        RECT 1064.990 52.330 1065.490 55.380 ;
        RECT 1069.960 52.240 1070.370 55.335 ;
        RECT 1069.000 50.580 1069.310 50.610 ;
        RECT 1059.800 46.860 1060.270 49.850 ;
        RECT 1062.150 43.875 1062.465 46.245 ;
        RECT 1063.770 45.920 1064.190 49.885 ;
        RECT 1060.435 41.165 1060.815 42.540 ;
        RECT 1062.875 40.135 1063.220 42.595 ;
        RECT 1064.510 41.815 1064.835 44.580 ;
        RECT 1065.495 43.850 1065.900 47.180 ;
        RECT 1069.000 44.480 1069.315 50.580 ;
        RECT 1070.145 40.875 1070.515 49.975 ;
        RECT 1071.090 41.940 1071.380 53.775 ;
        RECT 1074.540 52.215 1074.950 55.310 ;
        RECT 1078.995 51.670 1079.305 54.185 ;
        RECT 1083.245 53.370 1083.625 53.750 ;
        RECT 1085.375 53.370 1085.755 53.750 ;
        RECT 1071.985 44.435 1072.315 50.630 ;
        RECT 1074.890 43.905 1075.345 47.180 ;
        RECT 1077.250 45.920 1077.795 49.860 ;
        RECT 1081.305 46.860 1081.740 49.870 ;
        RECT 1076.445 41.815 1076.770 44.580 ;
        RECT 1078.960 43.910 1079.375 46.300 ;
        RECT 1082.500 42.485 1082.830 53.180 ;
        RECT 1083.935 46.820 1084.320 52.605 ;
        RECT 1080.690 41.080 1081.025 42.430 ;
        RECT 1084.295 42.065 1084.720 46.340 ;
        RECT 1085.995 43.830 1086.295 50.870 ;
        RECT 1087.115 43.225 1087.415 50.155 ;
        RECT 1088.425 43.825 1088.725 50.175 ;
        RECT 1082.955 41.155 1083.335 41.535 ;
        RECT 1085.150 41.140 1085.530 41.520 ;
        RECT 1089.020 41.080 1089.310 50.860 ;
        RECT 1089.740 43.855 1090.035 50.680 ;
        RECT 1090.870 43.315 1091.170 50.125 ;
        RECT 1091.660 43.910 1091.970 53.950 ;
        RECT 1100.850 52.195 1101.230 52.575 ;
        RECT 1092.455 43.840 1092.755 50.670 ;
        RECT 1093.580 43.225 1093.880 50.165 ;
        RECT 1095.030 43.100 1095.310 46.135 ;
        RECT 1095.790 43.800 1096.070 50.160 ;
        RECT 1096.640 43.800 1096.940 50.620 ;
        RECT 1097.780 43.055 1098.080 50.210 ;
        RECT 1098.425 47.245 1098.805 47.625 ;
        RECT 1098.425 45.190 1098.805 45.570 ;
        RECT 1100.275 45.070 1100.590 49.395 ;
        RECT 1100.885 47.145 1101.165 48.675 ;
        RECT 1101.455 43.830 1101.755 50.870 ;
        RECT 1102.575 43.225 1102.875 50.155 ;
        RECT 1103.230 44.585 1103.530 48.645 ;
        RECT 1103.885 43.825 1104.185 50.175 ;
        RECT 1100.750 42.020 1101.130 42.400 ;
        RECT 1104.480 41.615 1104.770 50.860 ;
        RECT 1105.200 43.855 1105.495 50.680 ;
        RECT 1106.330 43.315 1106.630 50.125 ;
        RECT 1107.120 43.910 1107.430 52.645 ;
        RECT 1107.915 43.840 1108.215 50.670 ;
        RECT 1109.040 43.225 1109.340 50.165 ;
        RECT 1109.720 44.570 1110.000 48.660 ;
        RECT 1110.490 43.100 1110.770 46.135 ;
        RECT 1111.250 43.800 1111.530 50.160 ;
        RECT 1112.100 43.800 1112.400 50.620 ;
        RECT 1113.240 43.055 1113.540 50.210 ;
        RECT 1115.580 48.825 1115.955 57.025 ;
        RECT 1117.325 48.020 1117.625 59.015 ;
        RECT 1118.275 47.095 1118.655 57.350 ;
        RECT 1119.145 44.940 1119.580 58.515 ;
        RECT 1174.855 57.675 1175.370 67.975 ;
        RECT 1176.540 56.570 1177.125 67.350 ;
        RECT 1178.035 64.825 1178.390 78.745 ;
        RECT 1241.380 78.115 1241.830 88.380 ;
        RECT 1179.660 65.730 1180.020 77.145 ;
        RECT 1242.545 76.575 1243.030 85.460 ;
        RECT 1249.210 76.310 1249.615 87.840 ;
        RECT 1251.285 78.210 1251.675 89.310 ;
        RECT 1254.710 81.690 1255.065 92.775 ;
        RECT 1256.035 86.545 1256.505 89.535 ;
        RECT 1256.670 80.850 1257.050 82.225 ;
        RECT 1257.440 81.670 1257.755 92.720 ;
        RECT 1258.455 91.415 1258.745 93.475 ;
        RECT 1261.225 92.015 1261.725 95.065 ;
        RECT 1266.195 91.925 1266.605 95.020 ;
        RECT 1265.235 90.265 1265.545 90.295 ;
        RECT 1258.385 83.560 1258.700 85.930 ;
        RECT 1260.005 85.605 1260.425 89.570 ;
        RECT 1259.110 79.820 1259.455 82.280 ;
        RECT 1260.745 81.500 1261.070 84.265 ;
        RECT 1261.730 83.535 1262.135 86.865 ;
        RECT 1265.235 84.165 1265.550 90.265 ;
        RECT 1266.380 80.560 1266.750 89.660 ;
        RECT 1267.325 81.625 1267.615 93.460 ;
        RECT 1270.775 91.900 1271.185 94.995 ;
        RECT 1275.230 91.355 1275.540 93.870 ;
        RECT 1279.480 93.055 1279.860 93.435 ;
        RECT 1281.610 93.055 1281.990 93.435 ;
        RECT 1268.220 84.120 1268.550 90.315 ;
        RECT 1271.125 83.590 1271.580 86.865 ;
        RECT 1273.485 85.605 1274.030 89.545 ;
        RECT 1272.680 81.500 1273.005 84.265 ;
        RECT 1275.195 83.595 1275.610 85.985 ;
        RECT 1276.225 82.155 1276.540 92.840 ;
        RECT 1277.540 86.545 1277.975 89.555 ;
        RECT 1278.735 82.170 1279.065 92.865 ;
        RECT 1279.415 87.915 1279.835 88.375 ;
        RECT 1280.170 86.505 1280.555 92.290 ;
        RECT 1280.915 87.910 1281.335 88.370 ;
        RECT 1279.550 85.025 1279.930 85.405 ;
        RECT 1276.925 80.765 1277.260 82.115 ;
        RECT 1280.530 81.750 1280.955 86.025 ;
        RECT 1281.615 85.000 1281.925 89.120 ;
        RECT 1282.230 83.515 1282.530 90.555 ;
        RECT 1283.350 82.910 1283.650 89.840 ;
        RECT 1284.005 84.270 1284.305 88.330 ;
        RECT 1284.660 83.510 1284.960 89.860 ;
        RECT 1279.190 80.840 1279.570 81.220 ;
        RECT 1281.385 80.825 1281.765 81.205 ;
        RECT 1285.255 80.765 1285.545 90.545 ;
        RECT 1285.975 83.540 1286.270 90.365 ;
        RECT 1287.105 83.000 1287.405 89.810 ;
        RECT 1287.895 83.595 1288.205 93.635 ;
        RECT 1288.690 83.525 1288.990 90.355 ;
        RECT 1289.815 82.910 1290.115 89.850 ;
        RECT 1290.495 84.255 1290.775 88.345 ;
        RECT 1291.265 82.785 1291.545 85.820 ;
        RECT 1292.025 83.485 1292.305 89.845 ;
        RECT 1292.875 83.485 1293.175 90.305 ;
        RECT 1294.015 82.740 1294.315 89.895 ;
        RECT 1294.685 88.695 1294.980 94.065 ;
        RECT 1295.260 87.865 1295.565 93.340 ;
        RECT 1297.085 91.880 1297.465 92.260 ;
        RECT 1294.660 86.930 1295.040 87.310 ;
        RECT 1294.660 84.875 1295.040 85.255 ;
        RECT 1296.510 84.755 1296.825 89.080 ;
        RECT 1297.120 86.830 1297.400 88.360 ;
        RECT 1297.690 83.515 1297.990 90.555 ;
        RECT 1299.465 84.270 1299.765 88.330 ;
        RECT 1296.985 81.705 1297.365 82.085 ;
        RECT 1300.715 81.300 1301.005 90.545 ;
        RECT 1302.565 83.000 1302.865 89.810 ;
        RECT 1303.355 83.595 1303.665 92.330 ;
        RECT 1304.150 83.525 1304.450 90.355 ;
        RECT 1305.955 84.255 1306.235 88.345 ;
        RECT 1306.725 82.785 1307.005 85.820 ;
        RECT 1309.475 82.740 1309.775 89.895 ;
        RECT 1311.760 88.600 1312.135 96.885 ;
        RECT 1313.505 87.880 1313.805 98.875 ;
        RECT 1183.445 68.960 1183.825 69.340 ;
        RECT 1183.435 68.210 1183.815 68.590 ;
        RECT 1183.480 67.525 1183.860 67.905 ;
        RECT 1183.445 66.855 1183.825 67.235 ;
        RECT 1184.160 63.780 1184.460 70.820 ;
        RECT 1185.280 63.175 1185.580 70.105 ;
        RECT 1185.935 64.535 1186.235 68.595 ;
        RECT 1186.590 63.775 1186.890 70.125 ;
        RECT 1187.185 65.650 1187.505 70.810 ;
        RECT 1187.905 63.805 1188.200 70.630 ;
        RECT 1189.035 63.265 1189.335 70.075 ;
        RECT 1189.825 63.860 1190.135 70.050 ;
        RECT 1190.620 63.790 1190.920 70.620 ;
        RECT 1191.745 63.175 1192.045 70.115 ;
        RECT 1192.425 64.520 1192.705 68.610 ;
        RECT 1193.195 63.050 1193.475 66.085 ;
        RECT 1193.955 63.750 1194.260 70.110 ;
        RECT 1194.805 63.750 1195.105 70.570 ;
        RECT 1195.945 63.005 1196.245 70.160 ;
        RECT 1196.610 68.960 1196.990 69.340 ;
        RECT 1198.880 68.960 1199.260 69.365 ;
        RECT 1196.615 68.210 1196.995 68.590 ;
        RECT 1198.885 68.210 1199.265 68.615 ;
        RECT 1196.615 67.195 1196.995 67.575 ;
        RECT 1198.400 65.775 1198.720 67.905 ;
        RECT 1196.830 62.485 1197.210 65.505 ;
        RECT 1199.010 64.935 1199.290 67.340 ;
        RECT 1199.620 63.780 1199.920 70.820 ;
        RECT 1200.740 63.175 1201.040 70.105 ;
        RECT 1201.395 64.535 1201.695 68.595 ;
        RECT 1202.050 63.775 1202.350 70.125 ;
        RECT 1202.645 65.650 1202.970 70.810 ;
        RECT 1203.365 63.805 1203.660 70.630 ;
        RECT 1204.495 63.265 1204.795 70.075 ;
        RECT 1205.285 63.860 1205.595 70.050 ;
        RECT 1206.080 63.790 1206.380 70.620 ;
        RECT 1207.205 63.175 1207.505 70.115 ;
        RECT 1207.885 64.520 1208.165 68.610 ;
        RECT 1208.655 63.050 1208.935 66.085 ;
        RECT 1209.415 63.750 1209.735 70.110 ;
        RECT 1210.265 63.750 1210.565 70.570 ;
        RECT 1211.405 63.005 1211.705 70.160 ;
        RECT 1212.345 68.960 1212.705 70.790 ;
        RECT 1212.040 65.150 1212.420 65.530 ;
        RECT 1212.745 61.035 1213.105 67.595 ;
        RECT 1213.885 65.785 1214.210 67.650 ;
        RECT 1214.525 67.440 1214.940 70.790 ;
        RECT 1214.550 62.440 1215.010 67.125 ;
        RECT 1215.335 64.985 1215.785 73.805 ;
        RECT 1216.195 62.610 1216.550 72.915 ;
        RECT 1216.860 68.215 1217.205 69.270 ;
        RECT 1217.520 66.810 1217.950 69.800 ;
        RECT 1215.265 61.095 1215.645 61.475 ;
        RECT 1218.155 61.115 1218.535 62.490 ;
        RECT 1218.925 61.935 1219.240 72.985 ;
        RECT 1219.940 71.680 1220.230 73.740 ;
        RECT 1222.725 72.280 1223.200 75.330 ;
        RECT 1227.680 72.190 1228.090 75.285 ;
        RECT 1226.720 70.530 1227.030 70.560 ;
        RECT 1219.860 63.825 1220.185 66.195 ;
        RECT 1221.510 65.870 1221.910 69.835 ;
        RECT 1220.595 60.085 1220.940 62.545 ;
        RECT 1222.230 61.765 1222.555 64.530 ;
        RECT 1223.215 63.800 1223.620 67.130 ;
        RECT 1226.720 64.430 1227.035 70.530 ;
        RECT 1227.865 60.825 1228.235 69.925 ;
        RECT 1228.810 61.890 1229.100 73.725 ;
        RECT 1232.260 72.165 1232.670 75.260 ;
        RECT 1236.715 71.620 1237.025 74.135 ;
        RECT 1229.705 64.385 1230.035 70.580 ;
        RECT 1232.625 63.855 1233.065 67.130 ;
        RECT 1235.005 65.870 1235.530 69.810 ;
        RECT 1234.165 61.765 1234.490 64.530 ;
        RECT 1236.680 63.860 1237.095 66.250 ;
        RECT 1237.710 62.420 1238.025 73.105 ;
        RECT 1239.040 66.810 1239.525 69.820 ;
        RECT 1240.220 62.435 1240.550 73.130 ;
        RECT 1238.410 61.030 1238.745 62.380 ;
        RECT 1150.055 42.130 1150.370 53.180 ;
        RECT 1153.890 52.475 1154.290 55.525 ;
        RECT 1158.810 52.385 1159.220 55.480 ;
        RECT 1163.390 52.360 1163.800 55.455 ;
        RECT 1151.725 40.280 1152.070 42.740 ;
        RECT 1168.840 42.615 1169.155 53.300 ;
        RECT 1174.025 45.405 1174.475 49.565 ;
        RECT 1175.725 48.385 1176.250 48.825 ;
        RECT 987.025 29.355 987.405 29.735 ;
        RECT 987.015 28.605 987.395 28.985 ;
        RECT 987.060 27.920 987.440 28.300 ;
        RECT 987.025 27.250 987.405 27.630 ;
        RECT 987.740 24.175 988.040 31.215 ;
        RECT 988.860 23.570 989.160 30.500 ;
        RECT 989.515 24.930 989.815 28.990 ;
        RECT 990.170 24.170 990.470 30.520 ;
        RECT 990.765 26.045 991.085 31.205 ;
        RECT 991.485 24.200 991.780 31.025 ;
        RECT 992.615 23.660 992.915 30.470 ;
        RECT 993.405 24.255 993.715 30.445 ;
        RECT 994.200 24.185 994.500 31.015 ;
        RECT 995.325 23.570 995.625 30.510 ;
        RECT 996.005 24.915 996.285 29.005 ;
        RECT 996.775 23.445 997.055 26.480 ;
        RECT 997.535 24.145 997.840 30.505 ;
        RECT 998.385 24.145 998.685 30.965 ;
        RECT 999.525 23.400 999.825 30.555 ;
        RECT 1000.190 29.355 1000.570 29.735 ;
        RECT 1002.460 29.355 1002.840 29.760 ;
        RECT 1000.195 28.605 1000.575 28.985 ;
        RECT 1002.465 28.605 1002.845 29.010 ;
        RECT 1000.195 27.590 1000.575 27.970 ;
        RECT 1001.980 26.170 1002.300 28.300 ;
        RECT 1000.410 22.880 1000.790 25.900 ;
        RECT 1002.590 25.330 1002.870 27.735 ;
        RECT 1003.200 24.175 1003.500 31.215 ;
        RECT 1004.320 23.570 1004.620 30.500 ;
        RECT 1004.975 24.930 1005.275 28.990 ;
        RECT 1005.630 24.170 1005.930 30.520 ;
        RECT 1006.225 26.045 1006.550 31.205 ;
        RECT 1006.945 24.200 1007.240 31.025 ;
        RECT 1008.075 23.660 1008.375 30.470 ;
        RECT 1008.865 24.255 1009.175 30.445 ;
        RECT 1009.660 24.185 1009.960 31.015 ;
        RECT 1010.785 23.570 1011.085 30.510 ;
        RECT 1011.465 24.915 1011.745 29.005 ;
        RECT 1012.235 23.445 1012.515 26.480 ;
        RECT 1012.995 24.145 1013.315 30.505 ;
        RECT 1013.845 24.145 1014.145 30.965 ;
        RECT 1014.985 23.400 1015.285 30.555 ;
        RECT 1015.925 29.355 1016.285 31.185 ;
        RECT 1015.620 25.545 1016.000 25.925 ;
        RECT 1016.325 21.430 1016.685 27.990 ;
        RECT 1017.465 26.180 1017.790 28.045 ;
        RECT 1018.105 27.835 1018.520 31.185 ;
        RECT 1018.130 22.835 1018.590 27.520 ;
        RECT 1018.915 25.380 1019.365 34.200 ;
        RECT 1019.775 23.005 1020.130 33.310 ;
        RECT 1020.440 28.610 1020.785 29.665 ;
        RECT 1021.100 27.205 1021.530 30.195 ;
        RECT 1018.845 21.490 1019.225 21.870 ;
        RECT 1021.735 21.510 1022.115 22.885 ;
        RECT 1022.505 22.330 1022.820 33.380 ;
        RECT 1023.520 32.075 1023.810 34.135 ;
        RECT 1026.305 32.675 1026.780 35.725 ;
        RECT 1031.260 32.585 1031.670 35.680 ;
        RECT 1030.300 30.925 1030.610 30.955 ;
        RECT 1023.440 24.220 1023.765 26.590 ;
        RECT 1025.090 26.265 1025.490 30.230 ;
        RECT 1024.175 20.480 1024.520 22.940 ;
        RECT 1025.810 22.160 1026.135 24.925 ;
        RECT 1026.795 24.195 1027.200 27.525 ;
        RECT 1030.300 24.825 1030.615 30.925 ;
        RECT 1031.445 21.220 1031.815 30.320 ;
        RECT 1032.390 22.285 1032.680 34.120 ;
        RECT 1035.840 32.560 1036.250 35.655 ;
        RECT 1040.295 32.015 1040.605 34.530 ;
        RECT 1033.285 24.780 1033.615 30.975 ;
        RECT 1036.205 24.250 1036.645 27.525 ;
        RECT 1038.585 26.265 1039.110 30.205 ;
        RECT 1037.745 22.160 1038.070 24.925 ;
        RECT 1040.260 24.255 1040.675 26.645 ;
        RECT 1041.290 22.815 1041.605 33.500 ;
        RECT 1042.620 27.205 1043.105 30.215 ;
        RECT 1043.800 22.830 1044.130 33.525 ;
        RECT 1049.080 29.125 1052.405 29.715 ;
        RECT 1049.080 28.510 1049.830 29.125 ;
        RECT 1050.985 25.670 1051.655 28.320 ;
        RECT 1041.990 21.425 1042.325 22.775 ;
        RECT 1052.945 9.515 1053.395 28.555 ;
        RECT 1054.735 8.740 1055.150 29.920 ;
        RECT 1058.475 22.340 1058.830 33.425 ;
        RECT 1062.220 32.065 1062.510 34.125 ;
        RECT 1064.990 32.665 1065.490 35.715 ;
        RECT 1069.960 32.575 1070.370 35.670 ;
        RECT 1069.000 30.915 1069.310 30.945 ;
        RECT 1059.800 27.195 1060.270 30.185 ;
        RECT 1062.150 24.210 1062.465 26.580 ;
        RECT 1063.770 26.255 1064.190 30.220 ;
        RECT 1060.435 21.500 1060.815 22.875 ;
        RECT 1062.875 20.470 1063.220 22.930 ;
        RECT 1064.510 22.150 1064.835 24.915 ;
        RECT 1065.495 24.185 1065.900 27.515 ;
        RECT 1069.000 24.815 1069.315 30.915 ;
        RECT 1070.145 21.210 1070.515 30.310 ;
        RECT 1071.090 22.275 1071.380 34.110 ;
        RECT 1074.540 32.550 1074.950 35.645 ;
        RECT 1078.995 32.005 1079.305 34.520 ;
        RECT 1083.245 33.705 1083.625 34.085 ;
        RECT 1085.375 33.705 1085.755 34.085 ;
        RECT 1071.985 24.770 1072.315 30.965 ;
        RECT 1074.890 24.240 1075.345 27.515 ;
        RECT 1077.250 26.255 1077.795 30.195 ;
        RECT 1081.305 27.195 1081.740 30.205 ;
        RECT 1076.445 22.150 1076.770 24.915 ;
        RECT 1078.960 24.245 1079.375 26.635 ;
        RECT 1082.500 22.820 1082.830 33.515 ;
        RECT 1083.935 27.155 1084.320 32.940 ;
        RECT 1080.690 21.415 1081.025 22.765 ;
        RECT 1084.295 22.400 1084.720 26.675 ;
        RECT 1085.995 24.165 1086.295 31.205 ;
        RECT 1087.115 23.560 1087.415 30.490 ;
        RECT 1088.425 24.160 1088.725 30.510 ;
        RECT 1082.955 21.490 1083.335 21.870 ;
        RECT 1085.150 21.475 1085.530 21.855 ;
        RECT 1089.020 21.415 1089.310 31.195 ;
        RECT 1089.740 24.190 1090.035 31.015 ;
        RECT 1090.870 23.650 1091.170 30.460 ;
        RECT 1091.660 24.245 1091.970 34.285 ;
        RECT 1100.850 32.530 1101.230 32.910 ;
        RECT 1092.455 24.175 1092.755 31.005 ;
        RECT 1093.580 23.560 1093.880 30.500 ;
        RECT 1095.030 23.435 1095.310 26.470 ;
        RECT 1095.790 24.135 1096.070 30.495 ;
        RECT 1096.640 24.135 1096.940 30.955 ;
        RECT 1097.780 23.390 1098.080 30.545 ;
        RECT 1098.425 27.580 1098.805 27.960 ;
        RECT 1098.425 25.525 1098.805 25.905 ;
        RECT 1100.275 25.405 1100.590 29.730 ;
        RECT 1100.885 27.480 1101.165 29.010 ;
        RECT 1101.455 24.165 1101.755 31.205 ;
        RECT 1102.575 23.560 1102.875 30.490 ;
        RECT 1103.230 24.920 1103.530 28.980 ;
        RECT 1103.885 24.160 1104.185 30.510 ;
        RECT 1100.750 22.355 1101.130 22.735 ;
        RECT 1104.480 21.950 1104.770 31.195 ;
        RECT 1105.200 24.190 1105.495 31.015 ;
        RECT 1106.330 23.650 1106.630 30.460 ;
        RECT 1107.120 24.245 1107.430 32.980 ;
        RECT 1107.915 24.175 1108.215 31.005 ;
        RECT 1109.040 23.560 1109.340 30.500 ;
        RECT 1109.720 24.905 1110.000 28.995 ;
        RECT 1110.490 23.435 1110.770 26.470 ;
        RECT 1111.250 24.135 1111.530 30.495 ;
        RECT 1112.100 24.135 1112.400 30.955 ;
        RECT 1113.240 23.390 1113.540 30.545 ;
        RECT 1115.165 29.310 1115.540 37.150 ;
        RECT 1117.020 28.560 1117.320 39.100 ;
        RECT 1118.275 27.435 1118.655 37.690 ;
        RECT 1119.145 25.280 1119.580 38.855 ;
        RECT 1174.855 38.120 1175.370 48.170 ;
        RECT 1176.540 36.765 1177.125 47.545 ;
        RECT 1178.130 45.060 1178.485 58.970 ;
        RECT 1241.475 58.340 1241.925 68.605 ;
        RECT 1179.755 45.980 1180.115 57.370 ;
        RECT 1242.640 56.800 1243.125 65.685 ;
        RECT 1249.470 56.155 1249.875 68.035 ;
        RECT 1251.545 58.055 1251.935 69.635 ;
        RECT 1254.815 61.975 1255.170 73.060 ;
        RECT 1256.140 66.830 1256.610 69.820 ;
        RECT 1256.775 61.135 1257.155 62.510 ;
        RECT 1257.545 61.955 1257.860 73.005 ;
        RECT 1258.560 71.700 1258.850 73.760 ;
        RECT 1261.330 72.300 1261.830 75.350 ;
        RECT 1266.300 72.210 1266.710 75.305 ;
        RECT 1265.340 70.550 1265.650 70.580 ;
        RECT 1258.490 63.845 1258.805 66.215 ;
        RECT 1260.110 65.890 1260.530 69.855 ;
        RECT 1259.215 60.105 1259.560 62.565 ;
        RECT 1260.850 61.785 1261.175 64.550 ;
        RECT 1261.835 63.820 1262.240 67.150 ;
        RECT 1265.340 64.450 1265.655 70.550 ;
        RECT 1266.485 60.845 1266.855 69.945 ;
        RECT 1267.430 61.910 1267.720 73.745 ;
        RECT 1270.880 72.185 1271.290 75.280 ;
        RECT 1275.335 71.640 1275.645 74.155 ;
        RECT 1279.585 73.340 1279.965 73.720 ;
        RECT 1281.715 73.340 1282.095 73.720 ;
        RECT 1268.325 64.405 1268.655 70.600 ;
        RECT 1271.230 63.875 1271.685 67.150 ;
        RECT 1273.590 65.890 1274.135 69.830 ;
        RECT 1272.785 61.785 1273.110 64.550 ;
        RECT 1275.300 63.880 1275.715 66.270 ;
        RECT 1276.330 62.440 1276.645 73.125 ;
        RECT 1277.645 66.830 1278.080 69.840 ;
        RECT 1278.840 62.455 1279.170 73.150 ;
        RECT 1279.520 68.200 1279.940 68.660 ;
        RECT 1280.275 66.790 1280.660 72.575 ;
        RECT 1281.020 68.195 1281.440 68.655 ;
        RECT 1279.655 65.310 1280.035 65.690 ;
        RECT 1277.030 61.050 1277.365 62.400 ;
        RECT 1280.635 62.035 1281.060 66.310 ;
        RECT 1281.720 65.285 1282.030 69.405 ;
        RECT 1282.335 63.800 1282.635 70.840 ;
        RECT 1283.455 63.195 1283.755 70.125 ;
        RECT 1284.110 64.555 1284.410 68.615 ;
        RECT 1284.765 63.795 1285.065 70.145 ;
        RECT 1279.295 61.125 1279.675 61.505 ;
        RECT 1281.490 61.110 1281.870 61.490 ;
        RECT 1285.360 61.050 1285.650 70.830 ;
        RECT 1286.080 63.825 1286.375 70.650 ;
        RECT 1287.210 63.285 1287.510 70.095 ;
        RECT 1288.000 63.880 1288.310 73.920 ;
        RECT 1288.795 63.810 1289.095 70.640 ;
        RECT 1289.920 63.195 1290.220 70.135 ;
        RECT 1290.600 64.540 1290.880 68.630 ;
        RECT 1291.370 63.070 1291.650 66.105 ;
        RECT 1292.130 63.770 1292.410 70.130 ;
        RECT 1292.980 63.770 1293.280 70.590 ;
        RECT 1294.120 63.025 1294.420 70.180 ;
        RECT 1294.790 68.980 1295.085 74.350 ;
        RECT 1295.365 68.150 1295.670 73.625 ;
        RECT 1297.190 72.165 1297.570 72.545 ;
        RECT 1294.765 67.215 1295.145 67.595 ;
        RECT 1294.765 65.160 1295.145 65.540 ;
        RECT 1296.615 65.040 1296.930 69.365 ;
        RECT 1297.225 67.115 1297.505 68.645 ;
        RECT 1297.795 63.800 1298.095 70.840 ;
        RECT 1299.570 64.555 1299.870 68.615 ;
        RECT 1297.090 61.990 1297.470 62.370 ;
        RECT 1300.820 61.585 1301.110 70.830 ;
        RECT 1302.670 63.285 1302.970 70.095 ;
        RECT 1303.460 63.880 1303.770 72.615 ;
        RECT 1304.255 63.810 1304.555 70.640 ;
        RECT 1306.060 64.540 1306.340 68.630 ;
        RECT 1306.830 63.070 1307.110 66.105 ;
        RECT 1309.580 63.025 1309.880 70.180 ;
        RECT 1311.660 68.900 1312.035 77.180 ;
        RECT 1313.405 68.060 1313.705 79.170 ;
        RECT 1183.395 49.150 1183.775 49.530 ;
        RECT 1183.385 48.400 1183.765 48.780 ;
        RECT 1183.430 47.715 1183.810 48.095 ;
        RECT 1183.395 47.045 1183.775 47.425 ;
        RECT 1184.110 43.970 1184.410 51.010 ;
        RECT 1185.230 43.365 1185.530 50.295 ;
        RECT 1185.885 44.725 1186.185 48.785 ;
        RECT 1186.540 43.965 1186.840 50.315 ;
        RECT 1187.135 45.840 1187.455 51.000 ;
        RECT 1187.855 43.995 1188.150 50.820 ;
        RECT 1188.985 43.455 1189.285 50.265 ;
        RECT 1189.775 44.050 1190.085 50.240 ;
        RECT 1190.570 43.980 1190.870 50.810 ;
        RECT 1191.695 43.365 1191.995 50.305 ;
        RECT 1192.375 44.710 1192.655 48.800 ;
        RECT 1193.145 43.240 1193.425 46.275 ;
        RECT 1193.905 43.940 1194.210 50.300 ;
        RECT 1194.755 43.940 1195.055 50.760 ;
        RECT 1195.895 43.195 1196.195 50.350 ;
        RECT 1196.560 49.150 1196.940 49.530 ;
        RECT 1198.830 49.150 1199.210 49.555 ;
        RECT 1196.565 48.400 1196.945 48.780 ;
        RECT 1198.835 48.400 1199.215 48.805 ;
        RECT 1196.565 47.385 1196.945 47.765 ;
        RECT 1198.350 45.965 1198.670 48.095 ;
        RECT 1196.780 42.675 1197.160 45.695 ;
        RECT 1198.960 45.125 1199.240 47.530 ;
        RECT 1199.570 43.970 1199.870 51.010 ;
        RECT 1200.690 43.365 1200.990 50.295 ;
        RECT 1201.345 44.725 1201.645 48.785 ;
        RECT 1202.000 43.965 1202.300 50.315 ;
        RECT 1202.595 45.840 1202.920 51.000 ;
        RECT 1203.315 43.995 1203.610 50.820 ;
        RECT 1204.445 43.455 1204.745 50.265 ;
        RECT 1205.235 44.050 1205.545 50.240 ;
        RECT 1206.030 43.980 1206.330 50.810 ;
        RECT 1207.155 43.365 1207.455 50.305 ;
        RECT 1207.835 44.710 1208.115 48.800 ;
        RECT 1208.605 43.240 1208.885 46.275 ;
        RECT 1209.365 43.940 1209.685 50.300 ;
        RECT 1210.215 43.940 1210.515 50.760 ;
        RECT 1211.355 43.195 1211.655 50.350 ;
        RECT 1212.295 49.150 1212.655 50.980 ;
        RECT 1211.990 45.340 1212.370 45.720 ;
        RECT 1212.695 41.225 1213.055 47.785 ;
        RECT 1213.835 45.975 1214.160 47.840 ;
        RECT 1214.475 47.630 1214.890 50.980 ;
        RECT 1214.500 42.630 1214.960 47.315 ;
        RECT 1215.285 45.175 1215.735 53.995 ;
        RECT 1216.145 42.800 1216.500 53.105 ;
        RECT 1216.810 48.405 1217.155 49.460 ;
        RECT 1217.470 47.000 1217.900 49.990 ;
        RECT 1215.215 41.285 1215.595 41.665 ;
        RECT 1218.105 41.305 1218.485 42.680 ;
        RECT 1218.875 42.125 1219.190 53.175 ;
        RECT 1219.890 51.870 1220.180 53.930 ;
        RECT 1222.675 52.470 1223.150 55.520 ;
        RECT 1227.630 52.380 1228.040 55.475 ;
        RECT 1226.670 50.720 1226.980 50.750 ;
        RECT 1219.810 44.015 1220.135 46.385 ;
        RECT 1221.460 46.060 1221.860 50.025 ;
        RECT 1220.545 40.275 1220.890 42.735 ;
        RECT 1222.180 41.955 1222.505 44.720 ;
        RECT 1223.165 43.990 1223.570 47.320 ;
        RECT 1226.670 44.620 1226.985 50.720 ;
        RECT 1227.815 41.015 1228.185 50.115 ;
        RECT 1228.760 42.080 1229.050 53.915 ;
        RECT 1232.210 52.355 1232.620 55.450 ;
        RECT 1236.665 51.810 1236.975 54.325 ;
        RECT 1229.655 44.575 1229.985 50.770 ;
        RECT 1232.575 44.045 1233.015 47.320 ;
        RECT 1234.955 46.060 1235.480 50.000 ;
        RECT 1234.115 41.955 1234.440 44.720 ;
        RECT 1236.630 44.050 1237.045 46.440 ;
        RECT 1237.660 42.610 1237.975 53.295 ;
        RECT 1238.990 47.000 1239.475 50.010 ;
        RECT 1240.170 42.625 1240.500 53.320 ;
        RECT 1238.360 41.220 1238.695 42.570 ;
        RECT 1150.030 22.400 1150.345 33.450 ;
        RECT 1153.865 32.745 1154.265 35.795 ;
        RECT 1158.785 32.655 1159.195 35.750 ;
        RECT 1163.365 32.630 1163.775 35.725 ;
        RECT 1151.700 20.550 1152.045 23.010 ;
        RECT 1168.815 22.885 1169.130 33.570 ;
        RECT 1174.050 25.600 1174.500 29.760 ;
        RECT 1175.750 28.580 1176.275 29.020 ;
        RECT 1058.495 3.825 1058.795 10.755 ;
        RECT 1059.150 5.185 1059.450 9.245 ;
        RECT 1059.805 4.425 1060.105 10.775 ;
        RECT 1061.120 4.455 1061.415 11.280 ;
        RECT 1064.960 3.825 1065.260 10.765 ;
        RECT 1065.640 5.170 1065.920 9.260 ;
        RECT 1067.170 4.400 1067.475 10.760 ;
        RECT 1068.020 4.400 1068.320 11.220 ;
        RECT 1069.750 7.840 1070.130 8.220 ;
        RECT 1069.760 5.795 1070.140 6.175 ;
        RECT 1174.850 5.440 1175.365 27.735 ;
        RECT 1176.535 7.655 1177.120 28.350 ;
        RECT 1178.130 25.220 1178.485 39.160 ;
        RECT 1241.475 38.530 1241.925 48.795 ;
        RECT 1179.755 26.010 1180.115 37.560 ;
        RECT 1242.640 36.990 1243.125 45.875 ;
        RECT 1249.580 36.265 1249.985 48.310 ;
        RECT 1251.655 38.165 1252.045 49.590 ;
        RECT 1254.815 42.005 1255.170 53.090 ;
        RECT 1256.140 46.860 1256.610 49.850 ;
        RECT 1256.775 41.165 1257.155 42.540 ;
        RECT 1257.545 41.985 1257.860 53.035 ;
        RECT 1258.560 51.730 1258.850 53.790 ;
        RECT 1261.330 52.330 1261.830 55.380 ;
        RECT 1266.300 52.240 1266.710 55.335 ;
        RECT 1265.340 50.580 1265.650 50.610 ;
        RECT 1258.490 43.875 1258.805 46.245 ;
        RECT 1260.110 45.920 1260.530 49.885 ;
        RECT 1259.215 40.135 1259.560 42.595 ;
        RECT 1260.850 41.815 1261.175 44.580 ;
        RECT 1261.835 43.850 1262.240 47.180 ;
        RECT 1265.340 44.480 1265.655 50.580 ;
        RECT 1266.485 40.875 1266.855 49.975 ;
        RECT 1267.430 41.940 1267.720 53.775 ;
        RECT 1270.880 52.215 1271.290 55.310 ;
        RECT 1275.335 51.670 1275.645 54.185 ;
        RECT 1279.585 53.370 1279.965 53.750 ;
        RECT 1281.715 53.370 1282.095 53.750 ;
        RECT 1268.325 44.435 1268.655 50.630 ;
        RECT 1271.230 43.905 1271.685 47.180 ;
        RECT 1273.590 45.920 1274.135 49.860 ;
        RECT 1272.785 41.815 1273.110 44.580 ;
        RECT 1275.300 43.910 1275.715 46.300 ;
        RECT 1276.330 42.470 1276.645 53.155 ;
        RECT 1277.645 46.860 1278.080 49.870 ;
        RECT 1278.840 42.485 1279.170 53.180 ;
        RECT 1279.520 48.230 1279.940 48.690 ;
        RECT 1280.275 46.820 1280.660 52.605 ;
        RECT 1281.020 48.225 1281.440 48.685 ;
        RECT 1279.655 45.340 1280.035 45.720 ;
        RECT 1277.030 41.080 1277.365 42.430 ;
        RECT 1280.635 42.065 1281.060 46.340 ;
        RECT 1281.720 45.315 1282.030 49.435 ;
        RECT 1282.335 43.830 1282.635 50.870 ;
        RECT 1283.455 43.225 1283.755 50.155 ;
        RECT 1284.110 44.585 1284.410 48.645 ;
        RECT 1284.765 43.825 1285.065 50.175 ;
        RECT 1279.295 41.155 1279.675 41.535 ;
        RECT 1281.490 41.140 1281.870 41.520 ;
        RECT 1285.360 41.080 1285.650 50.860 ;
        RECT 1286.080 43.855 1286.375 50.680 ;
        RECT 1287.210 43.315 1287.510 50.125 ;
        RECT 1288.000 43.910 1288.310 53.950 ;
        RECT 1288.795 43.840 1289.095 50.670 ;
        RECT 1289.920 43.225 1290.220 50.165 ;
        RECT 1290.600 44.570 1290.880 48.660 ;
        RECT 1291.370 43.100 1291.650 46.135 ;
        RECT 1292.130 43.800 1292.410 50.160 ;
        RECT 1292.980 43.800 1293.280 50.620 ;
        RECT 1294.120 43.055 1294.420 50.210 ;
        RECT 1294.790 49.010 1295.085 54.380 ;
        RECT 1295.365 48.180 1295.670 53.655 ;
        RECT 1297.190 52.195 1297.570 52.575 ;
        RECT 1294.765 47.245 1295.145 47.625 ;
        RECT 1294.765 45.190 1295.145 45.570 ;
        RECT 1296.615 45.070 1296.930 49.395 ;
        RECT 1297.225 47.145 1297.505 48.675 ;
        RECT 1297.795 43.830 1298.095 50.870 ;
        RECT 1299.570 44.585 1299.870 48.645 ;
        RECT 1297.090 42.020 1297.470 42.400 ;
        RECT 1300.820 41.615 1301.110 50.860 ;
        RECT 1302.670 43.315 1302.970 50.125 ;
        RECT 1303.460 43.910 1303.770 52.645 ;
        RECT 1304.255 43.840 1304.555 50.670 ;
        RECT 1306.060 44.570 1306.340 48.660 ;
        RECT 1306.830 43.100 1307.110 46.135 ;
        RECT 1309.580 43.055 1309.880 50.210 ;
        RECT 1311.920 48.825 1312.295 57.025 ;
        RECT 1313.665 48.020 1313.965 59.015 ;
        RECT 1183.365 29.355 1183.745 29.735 ;
        RECT 1183.355 28.605 1183.735 28.985 ;
        RECT 1183.400 27.920 1183.780 28.300 ;
        RECT 1183.365 27.250 1183.745 27.630 ;
        RECT 1184.080 24.175 1184.380 31.215 ;
        RECT 1185.200 23.570 1185.500 30.500 ;
        RECT 1185.855 24.930 1186.155 28.990 ;
        RECT 1186.510 24.170 1186.810 30.520 ;
        RECT 1187.105 26.045 1187.425 31.205 ;
        RECT 1187.825 24.200 1188.120 31.025 ;
        RECT 1188.955 23.660 1189.255 30.470 ;
        RECT 1189.745 24.255 1190.055 30.445 ;
        RECT 1190.540 24.185 1190.840 31.015 ;
        RECT 1191.665 23.570 1191.965 30.510 ;
        RECT 1192.345 24.915 1192.625 29.005 ;
        RECT 1193.115 23.445 1193.395 26.480 ;
        RECT 1193.875 24.145 1194.180 30.505 ;
        RECT 1194.725 24.145 1195.025 30.965 ;
        RECT 1195.865 23.400 1196.165 30.555 ;
        RECT 1196.530 29.355 1196.910 29.735 ;
        RECT 1198.800 29.355 1199.180 29.760 ;
        RECT 1196.535 28.605 1196.915 28.985 ;
        RECT 1198.805 28.605 1199.185 29.010 ;
        RECT 1196.535 27.590 1196.915 27.970 ;
        RECT 1198.320 26.170 1198.640 28.300 ;
        RECT 1196.750 22.880 1197.130 25.900 ;
        RECT 1198.930 25.330 1199.210 27.735 ;
        RECT 1199.540 24.175 1199.840 31.215 ;
        RECT 1200.660 23.570 1200.960 30.500 ;
        RECT 1201.315 24.930 1201.615 28.990 ;
        RECT 1201.970 24.170 1202.270 30.520 ;
        RECT 1202.565 26.045 1202.890 31.205 ;
        RECT 1203.285 24.200 1203.580 31.025 ;
        RECT 1204.415 23.660 1204.715 30.470 ;
        RECT 1205.205 24.255 1205.515 30.445 ;
        RECT 1206.000 24.185 1206.300 31.015 ;
        RECT 1207.125 23.570 1207.425 30.510 ;
        RECT 1207.805 24.915 1208.085 29.005 ;
        RECT 1208.575 23.445 1208.855 26.480 ;
        RECT 1209.335 24.145 1209.655 30.505 ;
        RECT 1210.185 24.145 1210.485 30.965 ;
        RECT 1211.325 23.400 1211.625 30.555 ;
        RECT 1212.265 29.355 1212.625 31.185 ;
        RECT 1211.960 25.545 1212.340 25.925 ;
        RECT 1212.665 21.430 1213.025 27.990 ;
        RECT 1213.805 26.180 1214.130 28.045 ;
        RECT 1214.445 27.835 1214.860 31.185 ;
        RECT 1214.470 22.835 1214.930 27.520 ;
        RECT 1215.255 25.380 1215.705 34.200 ;
        RECT 1216.115 23.005 1216.470 33.310 ;
        RECT 1216.780 28.610 1217.125 29.665 ;
        RECT 1217.440 27.205 1217.870 30.195 ;
        RECT 1215.185 21.490 1215.565 21.870 ;
        RECT 1218.075 21.510 1218.455 22.885 ;
        RECT 1218.845 22.330 1219.160 33.380 ;
        RECT 1219.860 32.075 1220.150 34.135 ;
        RECT 1222.645 32.675 1223.120 35.725 ;
        RECT 1227.600 32.585 1228.010 35.680 ;
        RECT 1226.640 30.925 1226.950 30.955 ;
        RECT 1219.780 24.220 1220.105 26.590 ;
        RECT 1221.430 26.265 1221.830 30.230 ;
        RECT 1220.515 20.480 1220.860 22.940 ;
        RECT 1222.150 22.160 1222.475 24.925 ;
        RECT 1223.135 24.195 1223.540 27.525 ;
        RECT 1226.640 24.825 1226.955 30.925 ;
        RECT 1227.785 21.220 1228.155 30.320 ;
        RECT 1228.730 22.285 1229.020 34.120 ;
        RECT 1232.180 32.560 1232.590 35.655 ;
        RECT 1236.635 32.015 1236.945 34.530 ;
        RECT 1229.625 24.780 1229.955 30.975 ;
        RECT 1232.545 24.250 1232.985 27.525 ;
        RECT 1234.925 26.265 1235.450 30.205 ;
        RECT 1234.085 22.160 1234.410 24.925 ;
        RECT 1236.600 24.255 1237.015 26.645 ;
        RECT 1237.630 22.815 1237.945 33.500 ;
        RECT 1238.960 27.205 1239.445 30.215 ;
        RECT 1240.140 22.830 1240.470 33.525 ;
        RECT 1245.420 29.125 1248.745 29.715 ;
        RECT 1245.420 28.510 1246.170 29.125 ;
        RECT 1247.325 25.670 1247.995 28.320 ;
        RECT 1238.330 21.425 1238.665 22.775 ;
        RECT 1249.285 9.515 1249.735 28.555 ;
        RECT 1251.075 8.740 1251.490 29.920 ;
        RECT 1254.815 22.340 1255.170 33.425 ;
        RECT 1256.140 27.195 1256.610 30.185 ;
        RECT 1256.775 21.500 1257.155 22.875 ;
        RECT 1257.545 22.320 1257.860 33.370 ;
        RECT 1258.560 32.065 1258.850 34.125 ;
        RECT 1261.330 32.665 1261.830 35.715 ;
        RECT 1266.300 32.575 1266.710 35.670 ;
        RECT 1265.340 30.915 1265.650 30.945 ;
        RECT 1258.490 24.210 1258.805 26.580 ;
        RECT 1260.110 26.255 1260.530 30.220 ;
        RECT 1259.215 20.470 1259.560 22.930 ;
        RECT 1260.850 22.150 1261.175 24.915 ;
        RECT 1261.835 24.185 1262.240 27.515 ;
        RECT 1265.340 24.815 1265.655 30.915 ;
        RECT 1266.485 21.210 1266.855 30.310 ;
        RECT 1267.430 22.275 1267.720 34.110 ;
        RECT 1270.880 32.550 1271.290 35.645 ;
        RECT 1275.335 32.005 1275.645 34.520 ;
        RECT 1279.585 33.705 1279.965 34.085 ;
        RECT 1281.715 33.705 1282.095 34.085 ;
        RECT 1268.325 24.770 1268.655 30.965 ;
        RECT 1271.230 24.240 1271.685 27.515 ;
        RECT 1273.590 26.255 1274.135 30.195 ;
        RECT 1272.785 22.150 1273.110 24.915 ;
        RECT 1275.300 24.245 1275.715 26.635 ;
        RECT 1276.330 22.805 1276.645 33.490 ;
        RECT 1277.645 27.195 1278.080 30.205 ;
        RECT 1278.840 22.820 1279.170 33.515 ;
        RECT 1279.520 28.565 1279.940 29.025 ;
        RECT 1280.275 27.155 1280.660 32.940 ;
        RECT 1281.020 28.560 1281.440 29.020 ;
        RECT 1279.655 25.675 1280.035 26.055 ;
        RECT 1277.030 21.415 1277.365 22.765 ;
        RECT 1280.635 22.400 1281.060 26.675 ;
        RECT 1281.720 25.650 1282.030 29.770 ;
        RECT 1282.335 24.165 1282.635 31.205 ;
        RECT 1283.455 23.560 1283.755 30.490 ;
        RECT 1284.110 24.920 1284.410 28.980 ;
        RECT 1284.765 24.160 1285.065 30.510 ;
        RECT 1279.295 21.490 1279.675 21.870 ;
        RECT 1281.490 21.475 1281.870 21.855 ;
        RECT 1285.360 21.415 1285.650 31.195 ;
        RECT 1286.080 24.190 1286.375 31.015 ;
        RECT 1287.210 23.650 1287.510 30.460 ;
        RECT 1288.000 24.245 1288.310 34.285 ;
        RECT 1288.795 24.175 1289.095 31.005 ;
        RECT 1289.920 23.560 1290.220 30.500 ;
        RECT 1290.600 24.905 1290.880 28.995 ;
        RECT 1291.370 23.435 1291.650 26.470 ;
        RECT 1292.130 24.135 1292.410 30.495 ;
        RECT 1292.980 24.135 1293.280 30.955 ;
        RECT 1294.120 23.390 1294.420 30.545 ;
        RECT 1294.790 29.345 1295.085 34.715 ;
        RECT 1295.365 28.515 1295.670 33.990 ;
        RECT 1297.190 32.530 1297.570 32.910 ;
        RECT 1294.765 27.580 1295.145 27.960 ;
        RECT 1294.765 25.525 1295.145 25.905 ;
        RECT 1296.615 25.405 1296.930 29.730 ;
        RECT 1297.225 27.480 1297.505 29.010 ;
        RECT 1297.795 24.165 1298.095 31.205 ;
        RECT 1299.570 24.920 1299.870 28.980 ;
        RECT 1297.090 22.355 1297.470 22.735 ;
        RECT 1300.820 21.950 1301.110 31.195 ;
        RECT 1302.670 23.650 1302.970 30.460 ;
        RECT 1303.460 24.245 1303.770 32.980 ;
        RECT 1304.255 24.175 1304.555 31.005 ;
        RECT 1306.060 24.905 1306.340 28.995 ;
        RECT 1306.830 23.435 1307.110 26.470 ;
        RECT 1309.580 23.390 1309.880 30.545 ;
        RECT 1311.505 29.310 1311.880 37.150 ;
        RECT 1313.360 28.560 1313.660 39.100 ;
        RECT 1255.490 5.185 1255.790 9.245 ;
        RECT 1261.980 5.170 1262.260 9.260 ;
      LAYER Metal3 ;
        RECT 1294.810 172.530 1310.830 172.940 ;
        RECT 101.400 171.960 103.995 172.390 ;
        RECT 297.765 171.960 300.360 172.390 ;
        RECT 494.165 171.910 496.760 172.340 ;
        RECT 690.540 171.945 693.135 172.375 ;
        RECT 886.880 171.945 889.475 172.375 ;
        RECT 1083.220 171.945 1085.815 172.375 ;
        RECT 1279.560 171.945 1282.155 172.375 ;
        RECT 1295.340 171.750 1310.820 172.205 ;
        RECT 102.080 170.835 119.450 171.175 ;
        RECT 298.445 170.835 315.815 171.175 ;
        RECT 494.845 170.785 512.215 171.125 ;
        RECT 691.220 170.820 708.590 171.160 ;
        RECT 887.560 170.820 904.930 171.160 ;
        RECT 1083.900 170.820 1101.270 171.160 ;
        RECT 1280.240 170.820 1297.610 171.160 ;
        RECT 34.180 169.130 36.885 169.470 ;
        RECT 230.545 169.130 233.250 169.470 ;
        RECT 426.945 169.080 429.650 169.420 ;
        RECT 623.320 169.115 626.025 169.455 ;
        RECT 819.660 169.115 822.365 169.455 ;
        RECT 1016.000 169.115 1018.705 169.455 ;
        RECT 1212.340 169.115 1215.045 169.455 ;
        RECT -0.230 168.020 5.750 168.030 ;
        RECT -4.025 167.725 5.750 168.020 ;
        RECT 18.445 167.715 21.190 168.045 ;
        RECT 192.145 167.735 202.115 168.030 ;
        RECT 196.135 167.725 202.115 167.735 ;
        RECT 214.810 167.715 217.555 168.045 ;
        RECT 584.855 168.015 589.085 168.035 ;
        RECT 388.535 167.980 392.765 167.990 ;
        RECT 388.535 167.695 398.515 167.980 ;
        RECT 392.535 167.675 398.515 167.695 ;
        RECT 411.210 167.665 413.955 167.995 ;
        RECT 584.855 167.740 594.890 168.015 ;
        RECT 588.910 167.710 594.890 167.740 ;
        RECT 607.585 167.700 610.330 168.030 ;
        RECT 781.220 168.015 785.450 168.040 ;
        RECT 781.220 167.745 791.230 168.015 ;
        RECT 785.250 167.710 791.230 167.745 ;
        RECT 803.925 167.700 806.670 168.030 ;
        RECT 977.605 168.015 981.835 168.025 ;
        RECT 977.605 167.730 987.570 168.015 ;
        RECT 981.590 167.710 987.570 167.730 ;
        RECT 1000.265 167.700 1003.010 168.030 ;
        RECT 1173.930 168.015 1178.160 168.030 ;
        RECT 1173.930 167.735 1183.910 168.015 ;
        RECT 1177.930 167.710 1183.910 167.735 ;
        RECT 1196.605 167.700 1199.350 168.030 ;
        RECT -2.130 167.285 0.185 167.345 ;
        RECT -2.130 167.000 5.730 167.285 ;
        RECT -0.215 166.990 5.730 167.000 ;
        RECT 18.450 166.965 21.190 167.295 ;
        RECT 194.040 167.285 196.355 167.355 ;
        RECT 194.040 167.010 202.095 167.285 ;
        RECT 196.150 166.990 202.095 167.010 ;
        RECT 214.815 166.965 217.555 167.295 ;
        RECT 390.430 167.235 392.745 167.315 ;
        RECT 586.750 167.270 589.065 167.360 ;
        RECT 390.430 166.970 398.495 167.235 ;
        RECT 392.550 166.940 398.495 166.970 ;
        RECT 411.215 166.915 413.955 167.245 ;
        RECT 586.750 167.015 594.870 167.270 ;
        RECT 588.925 166.975 594.870 167.015 ;
        RECT 607.590 166.950 610.330 167.280 ;
        RECT 783.115 167.270 785.430 167.365 ;
        RECT 783.115 167.020 791.210 167.270 ;
        RECT 785.265 166.975 791.210 167.020 ;
        RECT 803.930 166.950 806.670 167.280 ;
        RECT 979.500 167.270 981.815 167.350 ;
        RECT 979.500 167.005 987.550 167.270 ;
        RECT 981.605 166.975 987.550 167.005 ;
        RECT 1000.270 166.950 1003.010 167.280 ;
        RECT 1175.825 167.270 1178.140 167.355 ;
        RECT 1175.825 167.010 1183.890 167.270 ;
        RECT 1177.945 166.975 1183.890 167.010 ;
        RECT 1196.610 166.950 1199.350 167.280 ;
        RECT 1279.510 166.885 1281.535 167.270 ;
        RECT -55.800 166.275 5.765 166.570 ;
        RECT 192.995 166.275 202.130 166.570 ;
        RECT 18.455 165.945 36.180 166.265 ;
        RECT 214.820 165.945 232.545 166.265 ;
        RECT -55.080 165.645 5.720 165.940 ;
        RECT 193.115 165.645 202.085 165.940 ;
        RECT 312.970 165.865 315.815 166.245 ;
        RECT 389.395 166.225 398.530 166.520 ;
        RECT 585.770 166.260 594.905 166.555 ;
        RECT 782.110 166.260 791.245 166.555 ;
        RECT 978.450 166.260 987.585 166.555 ;
        RECT 1174.790 166.260 1183.925 166.555 ;
        RECT 411.220 165.895 428.945 166.215 ;
        RECT -55.080 165.635 0.070 165.645 ;
        RECT 389.515 165.595 398.485 165.890 ;
        RECT 509.370 165.815 512.215 166.195 ;
        RECT 607.595 165.930 625.320 166.250 ;
        RECT 585.890 165.630 594.860 165.925 ;
        RECT 705.745 165.850 708.590 166.230 ;
        RECT 803.935 165.930 821.660 166.250 ;
        RECT 782.230 165.630 791.200 165.925 ;
        RECT 902.085 165.850 904.930 166.230 ;
        RECT 1000.275 165.930 1018.000 166.250 ;
        RECT 978.570 165.630 987.540 165.925 ;
        RECT 1098.425 165.850 1101.270 166.230 ;
        RECT 1196.615 165.930 1214.340 166.250 ;
        RECT 1174.910 165.630 1183.880 165.925 ;
        RECT 1294.765 165.850 1297.610 166.230 ;
        RECT 196.155 164.570 217.040 164.865 ;
        RECT 392.555 164.520 413.440 164.815 ;
        RECT 588.930 164.555 609.815 164.850 ;
        RECT 785.270 164.555 806.155 164.850 ;
        RECT 981.610 164.555 1002.495 164.850 ;
        RECT 1177.950 164.555 1198.835 164.850 ;
        RECT 33.870 163.825 37.770 164.310 ;
        RECT 196.155 163.705 217.625 164.000 ;
        RECT 230.235 163.825 234.135 164.310 ;
        RECT 312.945 163.790 315.230 164.215 ;
        RECT 392.555 163.655 414.025 163.950 ;
        RECT 426.635 163.775 430.535 164.260 ;
        RECT 509.345 163.740 511.630 164.165 ;
        RECT 588.930 163.690 610.400 163.985 ;
        RECT 623.010 163.810 626.910 164.295 ;
        RECT 705.720 163.775 708.005 164.200 ;
        RECT 785.270 163.690 806.740 163.985 ;
        RECT 819.350 163.810 823.250 164.295 ;
        RECT 902.060 163.775 904.345 164.200 ;
        RECT 981.610 163.690 1003.080 163.985 ;
        RECT 1015.690 163.810 1019.590 164.295 ;
        RECT 1098.400 163.775 1100.685 164.200 ;
        RECT 1177.950 163.690 1199.420 163.985 ;
        RECT 1212.030 163.810 1215.930 164.295 ;
        RECT 1279.675 163.935 1282.155 164.335 ;
        RECT 1294.740 163.775 1297.025 164.200 ;
        RECT 18.620 161.170 36.920 161.555 ;
        RECT 214.985 161.170 233.285 161.555 ;
        RECT 411.385 161.120 429.685 161.505 ;
        RECT 607.760 161.155 626.060 161.540 ;
        RECT 804.100 161.155 822.400 161.540 ;
        RECT 1000.440 161.155 1018.740 161.540 ;
        RECT 1196.780 161.155 1215.080 161.540 ;
        RECT 102.335 160.635 119.520 161.120 ;
        RECT 298.700 160.635 315.885 161.120 ;
        RECT 495.100 160.585 512.285 161.070 ;
        RECT 691.475 160.620 708.660 161.105 ;
        RECT 887.815 160.620 905.000 161.105 ;
        RECT 1084.155 160.620 1101.340 161.105 ;
        RECT 1280.495 160.620 1297.680 161.105 ;
        RECT 34.500 159.850 37.565 160.175 ;
        RECT 101.145 159.720 103.740 160.170 ;
        RECT 230.865 159.850 233.930 160.175 ;
        RECT 297.510 159.720 300.105 160.170 ;
        RECT 427.265 159.800 430.330 160.125 ;
        RECT 493.910 159.670 496.505 160.120 ;
        RECT 623.640 159.835 626.705 160.160 ;
        RECT 690.285 159.705 692.880 160.155 ;
        RECT 819.980 159.835 823.045 160.160 ;
        RECT 886.625 159.705 889.220 160.155 ;
        RECT 1016.320 159.835 1019.385 160.160 ;
        RECT 1082.965 159.705 1085.560 160.155 ;
        RECT 1212.660 159.835 1215.725 160.160 ;
        RECT 1279.305 159.705 1281.900 160.155 ;
        RECT -0.070 157.095 63.810 157.515 ;
        RECT 72.485 157.220 135.930 157.840 ;
        RECT 137.185 156.775 193.955 157.270 ;
        RECT 196.295 157.095 260.175 157.515 ;
        RECT 268.850 157.220 332.295 157.840 ;
        RECT 333.575 156.735 390.345 157.230 ;
        RECT 392.695 157.045 456.575 157.465 ;
        RECT 465.250 157.170 528.695 157.790 ;
        RECT 529.895 156.780 586.665 157.275 ;
        RECT 589.070 157.080 652.950 157.500 ;
        RECT 661.625 157.205 725.070 157.825 ;
        RECT 726.260 156.785 783.030 157.280 ;
        RECT 785.410 157.080 849.290 157.500 ;
        RECT 857.965 157.205 921.410 157.825 ;
        RECT 922.645 156.770 979.415 157.265 ;
        RECT 981.750 157.080 1045.630 157.500 ;
        RECT 1054.305 157.205 1117.750 157.825 ;
        RECT 1118.970 156.775 1175.740 157.270 ;
        RECT 1178.090 157.080 1241.970 157.500 ;
        RECT 1250.645 157.205 1314.090 157.825 ;
        RECT 1.570 155.550 65.010 156.040 ;
        RECT 70.390 155.265 134.115 155.835 ;
        RECT 136.290 155.535 195.505 156.135 ;
        RECT 197.935 155.550 261.375 156.040 ;
        RECT 266.755 155.265 330.480 155.835 ;
        RECT 332.680 155.495 391.895 156.095 ;
        RECT 394.335 155.500 457.775 155.990 ;
        RECT 463.155 155.215 526.880 155.785 ;
        RECT 529.000 155.540 588.215 156.140 ;
        RECT 590.710 155.535 654.150 156.025 ;
        RECT 659.530 155.250 723.255 155.820 ;
        RECT 725.365 155.545 784.580 156.145 ;
        RECT 787.050 155.535 850.490 156.025 ;
        RECT 855.870 155.250 919.595 155.820 ;
        RECT 921.750 155.530 980.965 156.130 ;
        RECT 983.390 155.535 1046.830 156.025 ;
        RECT 1052.210 155.250 1115.935 155.820 ;
        RECT 1118.075 155.535 1177.290 156.135 ;
        RECT 1179.730 155.535 1243.170 156.025 ;
        RECT 1248.550 155.250 1312.275 155.820 ;
        RECT 1294.610 152.805 1310.630 153.215 ;
        RECT 101.200 152.235 103.795 152.665 ;
        RECT 297.565 152.235 300.160 152.665 ;
        RECT 493.965 152.185 496.560 152.615 ;
        RECT 690.340 152.220 692.935 152.650 ;
        RECT 886.680 152.220 889.275 152.650 ;
        RECT 1083.020 152.220 1085.615 152.650 ;
        RECT 1279.360 152.220 1281.955 152.650 ;
        RECT 1295.140 152.025 1310.620 152.480 ;
        RECT 101.880 151.110 119.250 151.450 ;
        RECT 298.245 151.110 315.615 151.450 ;
        RECT 494.645 151.060 512.015 151.400 ;
        RECT 691.020 151.095 708.390 151.435 ;
        RECT 887.360 151.095 904.730 151.435 ;
        RECT 1083.700 151.095 1101.070 151.435 ;
        RECT 1280.040 151.095 1297.410 151.435 ;
        RECT 34.135 149.440 36.840 149.780 ;
        RECT 230.500 149.440 233.205 149.780 ;
        RECT 426.900 149.390 429.605 149.730 ;
        RECT 623.275 149.425 625.980 149.765 ;
        RECT 819.615 149.425 822.320 149.765 ;
        RECT 1015.955 149.425 1018.660 149.765 ;
        RECT 1212.295 149.425 1215.000 149.765 ;
        RECT -0.275 148.305 5.705 148.340 ;
        RECT -4.110 148.035 5.705 148.305 ;
        RECT -4.110 148.010 0.120 148.035 ;
        RECT 18.400 148.025 21.145 148.355 ;
        RECT 196.090 148.315 202.070 148.340 ;
        RECT 192.060 148.035 202.070 148.315 ;
        RECT 192.060 148.020 196.290 148.035 ;
        RECT 214.765 148.025 217.510 148.355 ;
        RECT 588.865 148.320 594.845 148.325 ;
        RECT 392.490 148.275 398.470 148.290 ;
        RECT 388.450 147.985 398.470 148.275 ;
        RECT 388.450 147.980 392.680 147.985 ;
        RECT 411.165 147.975 413.910 148.305 ;
        RECT 584.770 148.025 594.845 148.320 ;
        RECT 588.865 148.020 594.845 148.025 ;
        RECT 607.540 148.010 610.285 148.340 ;
        RECT 781.135 148.030 791.185 148.325 ;
        RECT 785.205 148.020 791.185 148.030 ;
        RECT 803.880 148.010 806.625 148.340 ;
        RECT 981.545 148.310 987.525 148.325 ;
        RECT 977.520 148.020 987.525 148.310 ;
        RECT 977.520 148.015 981.750 148.020 ;
        RECT 1000.220 148.010 1002.965 148.340 ;
        RECT 1177.885 148.315 1183.865 148.325 ;
        RECT 1173.845 148.020 1183.865 148.315 ;
        RECT 1196.560 148.010 1199.305 148.340 ;
        RECT -2.235 147.595 0.100 147.630 ;
        RECT -2.235 147.300 5.685 147.595 ;
        RECT -2.235 147.285 0.100 147.300 ;
        RECT 18.405 147.275 21.145 147.605 ;
        RECT 193.935 147.595 196.270 147.640 ;
        RECT 193.935 147.300 202.050 147.595 ;
        RECT 193.935 147.295 196.270 147.300 ;
        RECT 214.770 147.275 217.510 147.605 ;
        RECT 390.325 147.545 392.660 147.600 ;
        RECT 586.645 147.580 588.980 147.645 ;
        RECT 390.325 147.255 398.450 147.545 ;
        RECT 392.505 147.250 398.450 147.255 ;
        RECT 411.170 147.225 413.910 147.555 ;
        RECT 586.645 147.300 594.825 147.580 ;
        RECT 588.880 147.285 594.825 147.300 ;
        RECT 607.545 147.260 610.285 147.590 ;
        RECT 783.010 147.580 785.345 147.650 ;
        RECT 783.010 147.305 791.165 147.580 ;
        RECT 785.220 147.285 791.165 147.305 ;
        RECT 803.885 147.260 806.625 147.590 ;
        RECT 979.395 147.580 981.730 147.635 ;
        RECT 979.395 147.290 987.505 147.580 ;
        RECT 981.560 147.285 987.505 147.290 ;
        RECT 1000.225 147.260 1002.965 147.590 ;
        RECT 1175.720 147.580 1178.055 147.640 ;
        RECT 1175.720 147.295 1183.845 147.580 ;
        RECT 1177.900 147.285 1183.845 147.295 ;
        RECT 1196.565 147.260 1199.305 147.590 ;
        RECT 1279.310 147.160 1281.335 147.545 ;
        RECT -3.415 146.855 5.720 146.880 ;
        RECT -55.920 146.585 5.720 146.855 ;
        RECT 192.950 146.585 202.085 146.880 ;
        RECT -55.920 146.560 0.035 146.585 ;
        RECT 18.410 146.255 36.135 146.575 ;
        RECT -3.295 146.225 5.675 146.250 ;
        RECT -55.130 145.955 5.675 146.225 ;
        RECT 116.405 146.140 119.250 146.520 ;
        RECT 214.775 146.255 232.500 146.575 ;
        RECT 389.350 146.535 398.485 146.830 ;
        RECT 585.725 146.570 594.860 146.865 ;
        RECT 782.065 146.570 791.200 146.865 ;
        RECT 978.405 146.570 987.540 146.865 ;
        RECT 1174.745 146.570 1183.880 146.865 ;
        RECT 193.070 145.955 202.040 146.250 ;
        RECT 312.770 146.140 315.615 146.520 ;
        RECT 411.175 146.205 428.900 146.525 ;
        RECT -55.130 145.920 -0.015 145.955 ;
        RECT 389.470 145.905 398.440 146.200 ;
        RECT 509.170 146.090 512.015 146.470 ;
        RECT 607.550 146.240 625.275 146.560 ;
        RECT 585.845 145.940 594.815 146.235 ;
        RECT 705.545 146.125 708.390 146.505 ;
        RECT 803.890 146.240 821.615 146.560 ;
        RECT 782.185 145.940 791.155 146.235 ;
        RECT 901.885 146.125 904.730 146.505 ;
        RECT 1000.230 146.240 1017.955 146.560 ;
        RECT 978.525 145.940 987.495 146.235 ;
        RECT 1098.225 146.125 1101.070 146.505 ;
        RECT 1196.570 146.240 1214.295 146.560 ;
        RECT 1174.865 145.940 1183.835 146.235 ;
        RECT 1294.565 146.125 1297.410 146.505 ;
        RECT -0.255 144.880 20.630 145.175 ;
        RECT 196.110 144.880 216.995 145.175 ;
        RECT 392.510 144.830 413.395 145.125 ;
        RECT 588.885 144.865 609.770 145.160 ;
        RECT 785.225 144.865 806.110 145.160 ;
        RECT 981.565 144.865 1002.450 145.160 ;
        RECT 1177.905 144.865 1198.790 145.160 ;
        RECT -0.255 144.015 21.215 144.310 ;
        RECT 33.825 144.135 37.725 144.620 ;
        RECT 116.380 144.065 118.665 144.490 ;
        RECT 196.110 144.015 217.580 144.310 ;
        RECT 230.190 144.135 234.090 144.620 ;
        RECT 312.745 144.065 315.030 144.490 ;
        RECT 392.510 143.965 413.980 144.260 ;
        RECT 426.590 144.085 430.490 144.570 ;
        RECT 509.145 144.015 511.430 144.440 ;
        RECT 588.885 144.000 610.355 144.295 ;
        RECT 622.965 144.120 626.865 144.605 ;
        RECT 705.520 144.050 707.805 144.475 ;
        RECT 785.225 144.000 806.695 144.295 ;
        RECT 819.305 144.120 823.205 144.605 ;
        RECT 901.860 144.050 904.145 144.475 ;
        RECT 981.565 144.000 1003.035 144.295 ;
        RECT 1015.645 144.120 1019.545 144.605 ;
        RECT 1098.200 144.050 1100.485 144.475 ;
        RECT 1177.905 144.000 1199.375 144.295 ;
        RECT 1211.985 144.120 1215.885 144.605 ;
        RECT 1279.475 144.210 1281.955 144.610 ;
        RECT 1294.540 144.050 1296.825 144.475 ;
        RECT 18.575 141.480 36.875 141.865 ;
        RECT 214.940 141.480 233.240 141.865 ;
        RECT 411.340 141.430 429.640 141.815 ;
        RECT 607.715 141.465 626.015 141.850 ;
        RECT 804.055 141.465 822.355 141.850 ;
        RECT 1000.395 141.465 1018.695 141.850 ;
        RECT 1196.735 141.465 1215.035 141.850 ;
        RECT 102.135 140.910 119.320 141.395 ;
        RECT 298.500 140.910 315.685 141.395 ;
        RECT 494.900 140.860 512.085 141.345 ;
        RECT 691.275 140.895 708.460 141.380 ;
        RECT 887.615 140.895 904.800 141.380 ;
        RECT 1083.955 140.895 1101.140 141.380 ;
        RECT 1280.295 140.895 1297.480 141.380 ;
        RECT 34.455 140.160 37.520 140.485 ;
        RECT 100.945 139.995 103.540 140.445 ;
        RECT 230.820 140.160 233.885 140.485 ;
        RECT 297.310 139.995 299.905 140.445 ;
        RECT 427.220 140.110 430.285 140.435 ;
        RECT 493.710 139.945 496.305 140.395 ;
        RECT 623.595 140.145 626.660 140.470 ;
        RECT 690.085 139.980 692.680 140.430 ;
        RECT 819.935 140.145 823.000 140.470 ;
        RECT 886.425 139.980 889.020 140.430 ;
        RECT 1016.275 140.145 1019.340 140.470 ;
        RECT 1082.765 139.980 1085.360 140.430 ;
        RECT 1212.615 140.145 1215.680 140.470 ;
        RECT 1279.105 139.980 1281.700 140.430 ;
        RECT -0.070 137.595 63.810 138.015 ;
        RECT 72.785 137.470 136.230 138.090 ;
        RECT 137.190 137.140 193.960 137.635 ;
        RECT 196.295 137.595 260.175 138.015 ;
        RECT 269.150 137.470 332.595 138.090 ;
        RECT 333.580 137.100 390.350 137.595 ;
        RECT 392.695 137.545 456.575 137.965 ;
        RECT 465.550 137.420 528.995 138.040 ;
        RECT 529.900 137.145 586.670 137.640 ;
        RECT 589.070 137.580 652.950 138.000 ;
        RECT 661.925 137.455 725.370 138.075 ;
        RECT 726.265 137.150 783.035 137.645 ;
        RECT 785.410 137.580 849.290 138.000 ;
        RECT 858.265 137.455 921.710 138.075 ;
        RECT 922.650 137.135 979.420 137.630 ;
        RECT 981.750 137.580 1045.630 138.000 ;
        RECT 1054.605 137.455 1118.050 138.075 ;
        RECT 1118.975 137.140 1175.745 137.635 ;
        RECT 1178.090 137.580 1241.970 138.000 ;
        RECT 1250.945 137.455 1314.390 138.075 ;
        RECT 1.570 136.050 65.010 136.540 ;
        RECT 70.690 135.515 134.415 136.085 ;
        RECT 136.295 135.900 195.510 136.500 ;
        RECT 197.935 136.050 261.375 136.540 ;
        RECT 267.055 135.515 330.780 136.085 ;
        RECT 332.685 135.860 391.900 136.460 ;
        RECT 394.335 136.000 457.775 136.490 ;
        RECT 463.455 135.465 527.180 136.035 ;
        RECT 529.005 135.905 588.220 136.505 ;
        RECT 590.710 136.035 654.150 136.525 ;
        RECT 659.830 135.500 723.555 136.070 ;
        RECT 725.370 135.910 784.585 136.510 ;
        RECT 787.050 136.035 850.490 136.525 ;
        RECT 856.170 135.500 919.895 136.070 ;
        RECT 921.755 135.895 980.970 136.495 ;
        RECT 983.390 136.035 1046.830 136.525 ;
        RECT 1052.510 135.500 1116.235 136.070 ;
        RECT 1118.080 135.900 1177.295 136.500 ;
        RECT 1179.730 136.035 1243.170 136.525 ;
        RECT 1248.850 135.500 1312.575 136.070 ;
        RECT 1294.765 133.160 1310.785 133.570 ;
        RECT 101.355 132.590 103.950 133.020 ;
        RECT 297.720 132.590 300.315 133.020 ;
        RECT 494.120 132.540 496.715 132.970 ;
        RECT 690.495 132.575 693.090 133.005 ;
        RECT 886.835 132.575 889.430 133.005 ;
        RECT 1083.175 132.575 1085.770 133.005 ;
        RECT 1279.515 132.575 1282.110 133.005 ;
        RECT 1295.295 132.380 1310.775 132.835 ;
        RECT 102.035 131.465 119.405 131.805 ;
        RECT 298.400 131.465 315.770 131.805 ;
        RECT 494.800 131.415 512.170 131.755 ;
        RECT 691.175 131.450 708.545 131.790 ;
        RECT 887.515 131.450 904.885 131.790 ;
        RECT 1083.855 131.450 1101.225 131.790 ;
        RECT 1280.195 131.450 1297.565 131.790 ;
        RECT 34.325 129.730 37.030 130.070 ;
        RECT 230.690 129.730 233.395 130.070 ;
        RECT 427.090 129.680 429.795 130.020 ;
        RECT 623.465 129.715 626.170 130.055 ;
        RECT 819.805 129.715 822.510 130.055 ;
        RECT 1016.145 129.715 1018.850 130.055 ;
        RECT 1212.485 129.715 1215.190 130.055 ;
        RECT -0.085 128.500 5.895 128.630 ;
        RECT -4.050 128.325 5.895 128.500 ;
        RECT -4.050 128.205 0.180 128.325 ;
        RECT 18.590 128.315 21.335 128.645 ;
        RECT 196.135 128.510 202.260 128.630 ;
        RECT 192.120 128.325 202.260 128.510 ;
        RECT 192.120 128.215 196.350 128.325 ;
        RECT 214.955 128.315 217.700 128.645 ;
        RECT 392.340 128.470 398.660 128.580 ;
        RECT 388.510 128.275 398.660 128.470 ;
        RECT 388.510 128.175 392.740 128.275 ;
        RECT 411.355 128.265 414.100 128.595 ;
        RECT 588.750 128.515 595.035 128.615 ;
        RECT 584.830 128.310 595.035 128.515 ;
        RECT 584.830 128.220 589.295 128.310 ;
        RECT 607.730 128.300 610.475 128.630 ;
        RECT 785.115 128.615 785.660 128.620 ;
        RECT 785.115 128.520 791.375 128.615 ;
        RECT 781.195 128.310 791.375 128.520 ;
        RECT 781.195 128.225 785.660 128.310 ;
        RECT 804.070 128.300 806.815 128.630 ;
        RECT 981.735 128.605 987.715 128.615 ;
        RECT 981.500 128.505 987.715 128.605 ;
        RECT 977.580 128.310 987.715 128.505 ;
        RECT 977.580 128.210 982.045 128.310 ;
        RECT 1000.410 128.300 1003.155 128.630 ;
        RECT 1178.075 128.610 1184.055 128.615 ;
        RECT 1177.825 128.510 1184.055 128.610 ;
        RECT 1173.905 128.310 1184.055 128.510 ;
        RECT 1173.905 128.215 1178.370 128.310 ;
        RECT 1196.750 128.300 1199.495 128.630 ;
        RECT -0.070 127.825 5.875 127.885 ;
        RECT -2.155 127.590 5.875 127.825 ;
        RECT -2.155 127.480 0.160 127.590 ;
        RECT 18.595 127.565 21.335 127.895 ;
        RECT 196.105 127.835 202.240 127.885 ;
        RECT 194.015 127.590 202.240 127.835 ;
        RECT 194.015 127.490 196.330 127.590 ;
        RECT 214.960 127.565 217.700 127.895 ;
        RECT 392.355 127.795 398.640 127.835 ;
        RECT 390.405 127.540 398.640 127.795 ;
        RECT 390.405 127.450 392.720 127.540 ;
        RECT 411.360 127.515 414.100 127.845 ;
        RECT 588.720 127.840 595.015 127.870 ;
        RECT 586.725 127.575 595.015 127.840 ;
        RECT 586.725 127.495 589.350 127.575 ;
        RECT 607.735 127.550 610.475 127.880 ;
        RECT 785.085 127.870 785.715 127.875 ;
        RECT 785.085 127.845 791.355 127.870 ;
        RECT 783.090 127.575 791.355 127.845 ;
        RECT 783.090 127.500 785.715 127.575 ;
        RECT 804.075 127.550 806.815 127.880 ;
        RECT 981.750 127.860 987.695 127.870 ;
        RECT 981.470 127.830 987.695 127.860 ;
        RECT 979.475 127.575 987.695 127.830 ;
        RECT 979.475 127.485 982.100 127.575 ;
        RECT 1000.415 127.550 1003.155 127.880 ;
        RECT 1178.090 127.865 1184.035 127.870 ;
        RECT 1177.795 127.835 1184.035 127.865 ;
        RECT 1175.800 127.575 1184.035 127.835 ;
        RECT 1175.800 127.490 1178.425 127.575 ;
        RECT 1196.755 127.550 1199.495 127.880 ;
        RECT 1279.465 127.515 1281.490 127.900 ;
        RECT -3.530 127.050 5.910 127.170 ;
        RECT -55.800 126.875 5.910 127.050 ;
        RECT 193.140 126.875 202.275 127.170 ;
        RECT -55.800 126.755 -3.310 126.875 ;
        RECT 18.600 126.545 36.325 126.865 ;
        RECT -3.105 126.420 5.865 126.540 ;
        RECT 116.560 126.495 119.405 126.875 ;
        RECT 214.965 126.545 232.690 126.865 ;
        RECT -55.090 126.245 5.865 126.420 ;
        RECT 193.260 126.245 202.230 126.540 ;
        RECT 312.925 126.495 315.770 126.875 ;
        RECT 389.540 126.825 398.675 127.120 ;
        RECT 585.915 126.860 595.050 127.155 ;
        RECT 782.255 126.860 791.390 127.155 ;
        RECT 978.595 126.860 987.730 127.155 ;
        RECT 1174.935 126.860 1184.070 127.155 ;
        RECT 411.365 126.495 429.090 126.815 ;
        RECT -55.090 126.115 0.045 126.245 ;
        RECT 389.660 126.195 398.630 126.490 ;
        RECT 509.325 126.445 512.170 126.825 ;
        RECT 607.740 126.530 625.465 126.850 ;
        RECT 586.035 126.230 595.005 126.525 ;
        RECT 705.700 126.480 708.545 126.860 ;
        RECT 804.080 126.530 821.805 126.850 ;
        RECT 782.375 126.230 791.345 126.525 ;
        RECT 902.040 126.480 904.885 126.860 ;
        RECT 1000.420 126.530 1018.145 126.850 ;
        RECT 978.715 126.230 987.685 126.525 ;
        RECT 1098.380 126.480 1101.225 126.860 ;
        RECT 1196.760 126.530 1214.485 126.850 ;
        RECT 1175.055 126.230 1184.025 126.525 ;
        RECT 1294.720 126.480 1297.565 126.860 ;
        RECT -0.065 125.170 20.820 125.465 ;
        RECT 196.300 125.170 217.185 125.465 ;
        RECT 392.700 125.120 413.585 125.415 ;
        RECT 589.075 125.155 609.960 125.450 ;
        RECT 785.415 125.155 806.300 125.450 ;
        RECT 981.755 125.155 1002.640 125.450 ;
        RECT 1178.095 125.155 1198.980 125.450 ;
        RECT -0.065 124.305 21.405 124.600 ;
        RECT 34.015 124.425 37.915 124.910 ;
        RECT 116.535 124.420 118.820 124.845 ;
        RECT 196.300 124.305 217.770 124.600 ;
        RECT 230.380 124.425 234.280 124.910 ;
        RECT 312.900 124.420 315.185 124.845 ;
        RECT 392.700 124.255 414.170 124.550 ;
        RECT 426.780 124.375 430.680 124.860 ;
        RECT 509.300 124.370 511.585 124.795 ;
        RECT 589.075 124.290 610.545 124.585 ;
        RECT 623.155 124.410 627.055 124.895 ;
        RECT 705.675 124.405 707.960 124.830 ;
        RECT 785.415 124.290 806.885 124.585 ;
        RECT 819.495 124.410 823.395 124.895 ;
        RECT 902.015 124.405 904.300 124.830 ;
        RECT 981.755 124.290 1003.225 124.585 ;
        RECT 1015.835 124.410 1019.735 124.895 ;
        RECT 1098.355 124.405 1100.640 124.830 ;
        RECT 1178.095 124.290 1199.565 124.585 ;
        RECT 1212.175 124.410 1216.075 124.895 ;
        RECT 1279.630 124.565 1282.110 124.965 ;
        RECT 1294.695 124.405 1296.980 124.830 ;
        RECT 18.765 121.770 37.065 122.155 ;
        RECT 215.130 121.770 233.430 122.155 ;
        RECT 102.290 121.265 119.475 121.750 ;
        RECT 298.655 121.265 315.840 121.750 ;
        RECT 411.530 121.720 429.830 122.105 ;
        RECT 607.905 121.755 626.205 122.140 ;
        RECT 804.245 121.755 822.545 122.140 ;
        RECT 1000.585 121.755 1018.885 122.140 ;
        RECT 1196.925 121.755 1215.225 122.140 ;
        RECT 495.055 121.215 512.240 121.700 ;
        RECT 691.430 121.250 708.615 121.735 ;
        RECT 887.770 121.250 904.955 121.735 ;
        RECT 1084.110 121.250 1101.295 121.735 ;
        RECT 1280.450 121.250 1297.635 121.735 ;
        RECT 34.645 120.450 37.710 120.775 ;
        RECT 101.100 120.350 103.695 120.800 ;
        RECT 231.010 120.450 234.075 120.775 ;
        RECT 297.465 120.350 300.060 120.800 ;
        RECT 427.410 120.400 430.475 120.725 ;
        RECT 493.865 120.300 496.460 120.750 ;
        RECT 623.785 120.435 626.850 120.760 ;
        RECT 690.240 120.335 692.835 120.785 ;
        RECT 820.125 120.435 823.190 120.760 ;
        RECT 886.580 120.335 889.175 120.785 ;
        RECT 1016.465 120.435 1019.530 120.760 ;
        RECT 1082.920 120.335 1085.515 120.785 ;
        RECT 1212.805 120.435 1215.870 120.760 ;
        RECT 1279.260 120.335 1281.855 120.785 ;
        RECT 0.140 117.555 64.020 117.975 ;
        RECT 72.805 117.810 136.250 118.430 ;
        RECT 137.190 117.375 193.960 117.870 ;
        RECT 196.505 117.555 260.385 117.975 ;
        RECT 269.170 117.810 332.615 118.430 ;
        RECT 333.580 117.335 390.350 117.830 ;
        RECT 392.905 117.505 456.785 117.925 ;
        RECT 465.570 117.760 529.015 118.380 ;
        RECT 529.900 117.380 586.670 117.875 ;
        RECT 589.280 117.540 653.160 117.960 ;
        RECT 661.945 117.795 725.390 118.415 ;
        RECT 726.265 117.385 783.035 117.880 ;
        RECT 785.620 117.540 849.500 117.960 ;
        RECT 858.285 117.795 921.730 118.415 ;
        RECT 922.650 117.370 979.420 117.865 ;
        RECT 981.960 117.540 1045.840 117.960 ;
        RECT 1054.625 117.795 1118.070 118.415 ;
        RECT 1118.975 117.375 1175.745 117.870 ;
        RECT 1178.300 117.540 1242.180 117.960 ;
        RECT 1250.965 117.795 1314.410 118.415 ;
        RECT 1.780 116.010 65.220 116.500 ;
        RECT 70.710 115.855 134.435 116.425 ;
        RECT 136.295 116.135 195.510 116.735 ;
        RECT 198.145 116.010 261.585 116.500 ;
        RECT 267.075 115.855 330.800 116.425 ;
        RECT 332.685 116.095 391.900 116.695 ;
        RECT 394.545 115.960 457.985 116.450 ;
        RECT 463.475 115.805 527.200 116.375 ;
        RECT 529.005 116.140 588.220 116.740 ;
        RECT 590.920 115.995 654.360 116.485 ;
        RECT 659.850 115.840 723.575 116.410 ;
        RECT 725.370 116.145 784.585 116.745 ;
        RECT 787.260 115.995 850.700 116.485 ;
        RECT 856.190 115.840 919.915 116.410 ;
        RECT 921.755 116.130 980.970 116.730 ;
        RECT 983.600 115.995 1047.040 116.485 ;
        RECT 1052.530 115.840 1116.255 116.410 ;
        RECT 1118.080 116.135 1177.295 116.735 ;
        RECT 1179.940 115.995 1243.380 116.485 ;
        RECT 1248.870 115.840 1312.595 116.410 ;
        RECT 1294.765 113.365 1310.785 113.775 ;
        RECT 101.355 112.795 103.950 113.225 ;
        RECT 297.720 112.795 300.315 113.225 ;
        RECT 494.120 112.745 496.715 113.175 ;
        RECT 690.495 112.780 693.090 113.210 ;
        RECT 886.835 112.780 889.430 113.210 ;
        RECT 1083.175 112.780 1085.770 113.210 ;
        RECT 1279.515 112.780 1282.110 113.210 ;
        RECT 1295.295 112.585 1310.775 113.040 ;
        RECT 102.035 111.670 119.405 112.010 ;
        RECT 298.400 111.670 315.770 112.010 ;
        RECT 494.800 111.620 512.170 111.960 ;
        RECT 691.175 111.655 708.545 111.995 ;
        RECT 887.515 111.655 904.885 111.995 ;
        RECT 1083.855 111.655 1101.225 111.995 ;
        RECT 1280.195 111.655 1297.565 111.995 ;
        RECT 34.130 109.890 36.835 110.230 ;
        RECT 230.495 109.890 233.200 110.230 ;
        RECT 426.895 109.840 429.600 110.180 ;
        RECT 623.270 109.875 625.975 110.215 ;
        RECT 819.610 109.875 822.315 110.215 ;
        RECT 1015.950 109.875 1018.655 110.215 ;
        RECT 1212.290 109.875 1214.995 110.215 ;
        RECT -0.280 108.730 5.700 108.790 ;
        RECT -4.120 108.485 5.700 108.730 ;
        RECT -4.120 108.435 0.110 108.485 ;
        RECT 18.395 108.475 21.140 108.805 ;
        RECT 196.085 108.740 202.065 108.790 ;
        RECT 192.050 108.485 202.065 108.740 ;
        RECT 192.050 108.445 196.280 108.485 ;
        RECT 214.760 108.475 217.505 108.805 ;
        RECT 392.485 108.700 398.465 108.740 ;
        RECT 388.440 108.435 398.465 108.700 ;
        RECT 388.440 108.405 392.670 108.435 ;
        RECT 411.160 108.425 413.905 108.755 ;
        RECT 588.860 108.745 594.840 108.775 ;
        RECT 584.760 108.470 594.840 108.745 ;
        RECT 584.760 108.450 588.990 108.470 ;
        RECT 607.535 108.460 610.280 108.790 ;
        RECT 785.200 108.750 791.180 108.775 ;
        RECT 781.125 108.470 791.180 108.750 ;
        RECT 781.125 108.455 785.355 108.470 ;
        RECT 803.875 108.460 806.620 108.790 ;
        RECT 981.540 108.735 987.520 108.775 ;
        RECT 977.510 108.470 987.520 108.735 ;
        RECT 977.510 108.440 981.740 108.470 ;
        RECT 1000.215 108.460 1002.960 108.790 ;
        RECT 1177.880 108.740 1183.860 108.775 ;
        RECT 1173.835 108.470 1183.860 108.740 ;
        RECT 1173.835 108.445 1178.065 108.470 ;
        RECT 1196.555 108.460 1199.300 108.790 ;
        RECT -2.225 108.045 0.090 108.055 ;
        RECT -2.225 107.750 5.680 108.045 ;
        RECT -2.225 107.710 0.090 107.750 ;
        RECT 18.400 107.725 21.140 108.055 ;
        RECT 193.945 108.045 196.260 108.065 ;
        RECT 193.945 107.750 202.045 108.045 ;
        RECT 193.945 107.720 196.260 107.750 ;
        RECT 214.765 107.725 217.505 108.055 ;
        RECT 586.655 108.030 588.970 108.070 ;
        RECT 390.335 107.995 392.650 108.025 ;
        RECT 390.335 107.700 398.445 107.995 ;
        RECT 390.335 107.680 392.650 107.700 ;
        RECT 411.165 107.675 413.905 108.005 ;
        RECT 586.655 107.735 594.820 108.030 ;
        RECT 586.655 107.725 588.970 107.735 ;
        RECT 607.540 107.710 610.280 108.040 ;
        RECT 783.020 108.030 785.335 108.075 ;
        RECT 783.020 107.735 791.160 108.030 ;
        RECT 783.020 107.730 785.335 107.735 ;
        RECT 803.880 107.710 806.620 108.040 ;
        RECT 979.405 108.030 981.720 108.060 ;
        RECT 979.405 107.735 987.500 108.030 ;
        RECT 979.405 107.715 981.720 107.735 ;
        RECT 1000.220 107.710 1002.960 108.040 ;
        RECT 1175.730 108.030 1178.045 108.065 ;
        RECT 1175.730 107.735 1183.840 108.030 ;
        RECT 1175.730 107.720 1178.045 107.735 ;
        RECT 1196.560 107.710 1199.300 108.040 ;
        RECT 1279.465 107.720 1281.490 108.105 ;
        RECT -3.420 107.280 5.715 107.330 ;
        RECT -55.865 107.035 5.715 107.280 ;
        RECT -55.865 106.985 0.025 107.035 ;
        RECT 18.405 106.705 36.130 107.025 ;
        RECT 116.560 106.700 119.405 107.080 ;
        RECT 192.945 107.035 202.080 107.330 ;
        RECT 214.770 106.705 232.495 107.025 ;
        RECT 312.925 106.700 315.770 107.080 ;
        RECT 389.345 106.985 398.480 107.280 ;
        RECT -3.300 106.650 5.670 106.700 ;
        RECT -55.140 106.405 5.670 106.650 ;
        RECT 193.065 106.405 202.035 106.700 ;
        RECT 411.170 106.655 428.895 106.975 ;
        RECT 509.325 106.650 512.170 107.030 ;
        RECT 585.720 107.020 594.855 107.315 ;
        RECT 607.545 106.690 625.270 107.010 ;
        RECT 705.700 106.685 708.545 107.065 ;
        RECT 782.060 107.020 791.195 107.315 ;
        RECT 803.885 106.690 821.610 107.010 ;
        RECT 902.040 106.685 904.885 107.065 ;
        RECT 978.400 107.020 987.535 107.315 ;
        RECT 1000.225 106.690 1017.950 107.010 ;
        RECT 1098.380 106.685 1101.225 107.065 ;
        RECT 1174.740 107.020 1183.875 107.315 ;
        RECT 1196.565 106.690 1214.290 107.010 ;
        RECT 1294.720 106.685 1297.565 107.065 ;
        RECT -55.140 106.345 -0.025 106.405 ;
        RECT 389.465 106.355 398.435 106.650 ;
        RECT 585.840 106.390 594.810 106.685 ;
        RECT 782.180 106.390 791.150 106.685 ;
        RECT 978.520 106.390 987.490 106.685 ;
        RECT 1174.860 106.390 1183.830 106.685 ;
        RECT -0.260 105.330 20.625 105.625 ;
        RECT 196.105 105.330 216.990 105.625 ;
        RECT 392.505 105.280 413.390 105.575 ;
        RECT 588.880 105.315 609.765 105.610 ;
        RECT 785.220 105.315 806.105 105.610 ;
        RECT 981.560 105.315 1002.445 105.610 ;
        RECT 1177.900 105.315 1198.785 105.610 ;
        RECT -0.260 104.465 21.210 104.760 ;
        RECT 33.820 104.585 37.720 105.070 ;
        RECT 116.535 104.625 118.820 105.050 ;
        RECT 196.105 104.465 217.575 104.760 ;
        RECT 230.185 104.585 234.085 105.070 ;
        RECT 312.900 104.625 315.185 105.050 ;
        RECT 392.505 104.415 413.975 104.710 ;
        RECT 426.585 104.535 430.485 105.020 ;
        RECT 509.300 104.575 511.585 105.000 ;
        RECT 588.880 104.450 610.350 104.745 ;
        RECT 622.960 104.570 626.860 105.055 ;
        RECT 705.675 104.610 707.960 105.035 ;
        RECT 785.220 104.450 806.690 104.745 ;
        RECT 819.300 104.570 823.200 105.055 ;
        RECT 902.015 104.610 904.300 105.035 ;
        RECT 981.560 104.450 1003.030 104.745 ;
        RECT 1015.640 104.570 1019.540 105.055 ;
        RECT 1098.355 104.610 1100.640 105.035 ;
        RECT 1177.900 104.450 1199.370 104.745 ;
        RECT 1211.980 104.570 1215.880 105.055 ;
        RECT 1279.630 104.770 1282.110 105.170 ;
        RECT 1294.695 104.610 1296.980 105.035 ;
        RECT 18.570 101.930 36.870 102.315 ;
        RECT 102.290 101.470 119.475 101.955 ;
        RECT 214.935 101.930 233.235 102.315 ;
        RECT 298.655 101.470 315.840 101.955 ;
        RECT 411.335 101.880 429.635 102.265 ;
        RECT 607.710 101.915 626.010 102.300 ;
        RECT 495.055 101.420 512.240 101.905 ;
        RECT 691.430 101.455 708.615 101.940 ;
        RECT 804.050 101.915 822.350 102.300 ;
        RECT 887.770 101.455 904.955 101.940 ;
        RECT 1000.390 101.915 1018.690 102.300 ;
        RECT 1084.110 101.455 1101.295 101.940 ;
        RECT 1196.730 101.915 1215.030 102.300 ;
        RECT 1280.450 101.455 1297.635 101.940 ;
        RECT 34.450 100.610 37.515 100.935 ;
        RECT 101.100 100.555 103.695 101.005 ;
        RECT 230.815 100.610 233.880 100.935 ;
        RECT 297.465 100.555 300.060 101.005 ;
        RECT 427.215 100.560 430.280 100.885 ;
        RECT 493.865 100.505 496.460 100.955 ;
        RECT 623.590 100.595 626.655 100.920 ;
        RECT 690.240 100.540 692.835 100.990 ;
        RECT 819.930 100.595 822.995 100.920 ;
        RECT 886.580 100.540 889.175 100.990 ;
        RECT 1016.270 100.595 1019.335 100.920 ;
        RECT 1082.920 100.540 1085.515 100.990 ;
        RECT 1212.610 100.595 1215.675 100.920 ;
        RECT 1279.260 100.540 1281.855 100.990 ;
        RECT 0.095 97.765 63.975 98.185 ;
        RECT 72.805 98.075 136.250 98.695 ;
        RECT 137.190 97.565 193.960 98.060 ;
        RECT 196.460 97.765 260.340 98.185 ;
        RECT 269.170 98.075 332.615 98.695 ;
        RECT 333.580 97.525 390.350 98.020 ;
        RECT 392.860 97.715 456.740 98.135 ;
        RECT 465.570 98.025 529.015 98.645 ;
        RECT 529.900 97.570 586.670 98.065 ;
        RECT 589.235 97.750 653.115 98.170 ;
        RECT 661.945 98.060 725.390 98.680 ;
        RECT 726.265 97.575 783.035 98.070 ;
        RECT 785.575 97.750 849.455 98.170 ;
        RECT 858.285 98.060 921.730 98.680 ;
        RECT 922.650 97.560 979.420 98.055 ;
        RECT 981.915 97.750 1045.795 98.170 ;
        RECT 1054.625 98.060 1118.070 98.680 ;
        RECT 1118.975 97.565 1175.745 98.060 ;
        RECT 1178.255 97.750 1242.135 98.170 ;
        RECT 1250.965 98.060 1314.410 98.680 ;
        RECT 1.735 96.220 65.175 96.710 ;
        RECT 70.710 96.120 134.435 96.690 ;
        RECT 136.295 96.325 195.510 96.925 ;
        RECT 198.100 96.220 261.540 96.710 ;
        RECT 267.075 96.120 330.800 96.690 ;
        RECT 332.685 96.285 391.900 96.885 ;
        RECT 394.500 96.170 457.940 96.660 ;
        RECT 463.475 96.070 527.200 96.640 ;
        RECT 529.005 96.330 588.220 96.930 ;
        RECT 590.875 96.205 654.315 96.695 ;
        RECT 659.850 96.105 723.575 96.675 ;
        RECT 725.370 96.335 784.585 96.935 ;
        RECT 787.215 96.205 850.655 96.695 ;
        RECT 856.190 96.105 919.915 96.675 ;
        RECT 921.755 96.320 980.970 96.920 ;
        RECT 983.555 96.205 1046.995 96.695 ;
        RECT 1052.530 96.105 1116.255 96.675 ;
        RECT 1118.080 96.325 1177.295 96.925 ;
        RECT 1179.895 96.205 1243.335 96.695 ;
        RECT 1248.870 96.105 1312.595 96.675 ;
        RECT 1294.685 93.610 1310.705 94.020 ;
        RECT 101.275 93.040 103.870 93.470 ;
        RECT 297.640 93.040 300.235 93.470 ;
        RECT 494.040 92.990 496.635 93.420 ;
        RECT 690.415 93.025 693.010 93.455 ;
        RECT 886.755 93.025 889.350 93.455 ;
        RECT 1083.095 93.025 1085.690 93.455 ;
        RECT 1279.435 93.025 1282.030 93.455 ;
        RECT 1295.215 92.830 1310.695 93.285 ;
        RECT 101.955 91.915 119.325 92.255 ;
        RECT 298.320 91.915 315.690 92.255 ;
        RECT 494.720 91.865 512.090 92.205 ;
        RECT 691.095 91.900 708.465 92.240 ;
        RECT 887.435 91.900 904.805 92.240 ;
        RECT 1083.775 91.900 1101.145 92.240 ;
        RECT 1280.115 91.900 1297.485 92.240 ;
        RECT 34.000 90.180 36.705 90.520 ;
        RECT 230.365 90.180 233.070 90.520 ;
        RECT 426.765 90.130 429.470 90.470 ;
        RECT 623.140 90.165 625.845 90.505 ;
        RECT 819.480 90.165 822.185 90.505 ;
        RECT 1015.820 90.165 1018.525 90.505 ;
        RECT 1212.160 90.165 1214.865 90.505 ;
        RECT -0.410 89.005 5.570 89.080 ;
        RECT -4.090 88.775 5.570 89.005 ;
        RECT -4.090 88.710 0.140 88.775 ;
        RECT 18.265 88.765 21.010 89.095 ;
        RECT 195.955 89.015 201.935 89.080 ;
        RECT 192.080 88.775 201.935 89.015 ;
        RECT 192.080 88.720 196.310 88.775 ;
        RECT 214.630 88.765 217.375 89.095 ;
        RECT 392.355 88.975 398.335 89.030 ;
        RECT 388.470 88.725 398.335 88.975 ;
        RECT 388.470 88.680 392.700 88.725 ;
        RECT 411.030 88.715 413.775 89.045 ;
        RECT 588.730 89.020 594.710 89.065 ;
        RECT 584.790 88.760 594.710 89.020 ;
        RECT 584.790 88.725 589.020 88.760 ;
        RECT 607.405 88.750 610.150 89.080 ;
        RECT 785.070 89.025 791.050 89.065 ;
        RECT 781.155 88.760 791.050 89.025 ;
        RECT 781.155 88.730 785.385 88.760 ;
        RECT 803.745 88.750 806.490 89.080 ;
        RECT 981.410 89.010 987.390 89.065 ;
        RECT 977.540 88.760 987.390 89.010 ;
        RECT 977.540 88.715 981.770 88.760 ;
        RECT 1000.085 88.750 1002.830 89.080 ;
        RECT 1177.750 89.015 1183.730 89.065 ;
        RECT 1173.865 88.760 1183.730 89.015 ;
        RECT 1173.865 88.720 1178.095 88.760 ;
        RECT 1196.425 88.750 1199.170 89.080 ;
        RECT -0.395 88.330 5.550 88.335 ;
        RECT -2.195 88.040 5.550 88.330 ;
        RECT -2.195 87.985 0.120 88.040 ;
        RECT 18.270 88.015 21.010 88.345 ;
        RECT 193.975 88.335 196.290 88.340 ;
        RECT 193.975 88.040 201.915 88.335 ;
        RECT 193.975 87.995 196.290 88.040 ;
        RECT 214.635 88.015 217.375 88.345 ;
        RECT 586.685 88.320 589.000 88.345 ;
        RECT 390.365 88.285 392.680 88.300 ;
        RECT 390.365 87.990 398.315 88.285 ;
        RECT 390.365 87.955 392.680 87.990 ;
        RECT 411.035 87.965 413.775 88.295 ;
        RECT 586.685 88.025 594.690 88.320 ;
        RECT 586.685 88.000 589.000 88.025 ;
        RECT 607.410 88.000 610.150 88.330 ;
        RECT 783.050 88.320 785.365 88.350 ;
        RECT 783.050 88.025 791.030 88.320 ;
        RECT 783.050 88.005 785.365 88.025 ;
        RECT 803.750 88.000 806.490 88.330 ;
        RECT 979.435 88.320 981.750 88.335 ;
        RECT 979.435 88.025 987.370 88.320 ;
        RECT 979.435 87.990 981.750 88.025 ;
        RECT 1000.090 88.000 1002.830 88.330 ;
        RECT 1175.760 88.320 1178.075 88.340 ;
        RECT 1175.760 88.025 1183.710 88.320 ;
        RECT 1175.760 87.995 1178.075 88.025 ;
        RECT 1196.430 88.000 1199.170 88.330 ;
        RECT 1279.385 87.965 1281.410 88.350 ;
        RECT -3.815 87.555 5.585 87.620 ;
        RECT -55.865 87.325 5.585 87.555 ;
        RECT 192.815 87.325 201.950 87.620 ;
        RECT -55.865 87.260 -3.525 87.325 ;
        RECT 18.275 86.995 36.000 87.315 ;
        RECT -3.430 86.925 5.540 86.990 ;
        RECT 116.480 86.945 119.325 87.325 ;
        RECT 214.640 86.995 232.365 87.315 ;
        RECT -55.150 86.695 5.540 86.925 ;
        RECT 192.935 86.695 201.905 86.990 ;
        RECT 312.845 86.945 315.690 87.325 ;
        RECT 389.215 87.275 398.350 87.570 ;
        RECT 585.590 87.310 594.725 87.605 ;
        RECT 781.930 87.310 791.065 87.605 ;
        RECT 978.270 87.310 987.405 87.605 ;
        RECT 1174.610 87.310 1183.745 87.605 ;
        RECT 411.040 86.945 428.765 87.265 ;
        RECT -55.150 86.620 0.005 86.695 ;
        RECT 389.335 86.645 398.305 86.940 ;
        RECT 509.245 86.895 512.090 87.275 ;
        RECT 607.415 86.980 625.140 87.300 ;
        RECT 585.710 86.680 594.680 86.975 ;
        RECT 705.620 86.930 708.465 87.310 ;
        RECT 803.755 86.980 821.480 87.300 ;
        RECT 782.050 86.680 791.020 86.975 ;
        RECT 901.960 86.930 904.805 87.310 ;
        RECT 1000.095 86.980 1017.820 87.300 ;
        RECT 978.390 86.680 987.360 86.975 ;
        RECT 1098.300 86.930 1101.145 87.310 ;
        RECT 1196.435 86.980 1214.160 87.300 ;
        RECT 1174.730 86.680 1183.700 86.975 ;
        RECT 1294.640 86.930 1297.485 87.310 ;
        RECT -0.390 85.620 20.495 85.915 ;
        RECT 195.975 85.620 216.860 85.915 ;
        RECT 392.375 85.570 413.260 85.865 ;
        RECT 588.750 85.605 609.635 85.900 ;
        RECT 785.090 85.605 805.975 85.900 ;
        RECT 981.430 85.605 1002.315 85.900 ;
        RECT 1177.770 85.605 1198.655 85.900 ;
        RECT -0.390 84.755 21.080 85.050 ;
        RECT 33.690 84.875 37.590 85.360 ;
        RECT 116.455 84.870 118.740 85.295 ;
        RECT 195.975 84.755 217.445 85.050 ;
        RECT 230.055 84.875 233.955 85.360 ;
        RECT 312.820 84.870 315.105 85.295 ;
        RECT 392.375 84.705 413.845 85.000 ;
        RECT 426.455 84.825 430.355 85.310 ;
        RECT 509.220 84.820 511.505 85.245 ;
        RECT 588.750 84.740 610.220 85.035 ;
        RECT 622.830 84.860 626.730 85.345 ;
        RECT 705.595 84.855 707.880 85.280 ;
        RECT 785.090 84.740 806.560 85.035 ;
        RECT 819.170 84.860 823.070 85.345 ;
        RECT 901.935 84.855 904.220 85.280 ;
        RECT 981.430 84.740 1002.900 85.035 ;
        RECT 1015.510 84.860 1019.410 85.345 ;
        RECT 1098.275 84.855 1100.560 85.280 ;
        RECT 1177.770 84.740 1199.240 85.035 ;
        RECT 1211.850 84.860 1215.750 85.345 ;
        RECT 1279.550 85.015 1282.030 85.415 ;
        RECT 1294.615 84.855 1296.900 85.280 ;
        RECT 18.440 82.220 36.740 82.605 ;
        RECT 214.805 82.220 233.105 82.605 ;
        RECT 102.210 81.715 119.395 82.200 ;
        RECT 298.575 81.715 315.760 82.200 ;
        RECT 411.205 82.170 429.505 82.555 ;
        RECT 607.580 82.205 625.880 82.590 ;
        RECT 803.920 82.205 822.220 82.590 ;
        RECT 1000.260 82.205 1018.560 82.590 ;
        RECT 1196.600 82.205 1214.900 82.590 ;
        RECT 494.975 81.665 512.160 82.150 ;
        RECT 691.350 81.700 708.535 82.185 ;
        RECT 887.690 81.700 904.875 82.185 ;
        RECT 1084.030 81.700 1101.215 82.185 ;
        RECT 1280.370 81.700 1297.555 82.185 ;
        RECT 34.320 80.900 37.385 81.225 ;
        RECT 101.020 80.800 103.615 81.250 ;
        RECT 230.685 80.900 233.750 81.225 ;
        RECT 297.385 80.800 299.980 81.250 ;
        RECT 427.085 80.850 430.150 81.175 ;
        RECT 493.785 80.750 496.380 81.200 ;
        RECT 623.460 80.885 626.525 81.210 ;
        RECT 690.160 80.785 692.755 81.235 ;
        RECT 819.800 80.885 822.865 81.210 ;
        RECT 886.500 80.785 889.095 81.235 ;
        RECT 1016.140 80.885 1019.205 81.210 ;
        RECT 1082.840 80.785 1085.435 81.235 ;
        RECT 1212.480 80.885 1215.545 81.210 ;
        RECT 1279.180 80.785 1281.775 81.235 ;
        RECT -0.210 78.135 63.670 78.555 ;
        RECT 72.705 78.370 136.150 78.990 ;
        RECT 137.180 77.915 193.950 78.410 ;
        RECT 196.155 78.135 260.035 78.555 ;
        RECT 269.070 78.370 332.515 78.990 ;
        RECT 333.570 77.875 390.340 78.370 ;
        RECT 392.555 78.085 456.435 78.505 ;
        RECT 465.470 78.320 528.915 78.940 ;
        RECT 529.890 77.920 586.660 78.415 ;
        RECT 588.930 78.120 652.810 78.540 ;
        RECT 661.845 78.355 725.290 78.975 ;
        RECT 726.255 77.925 783.025 78.420 ;
        RECT 785.270 78.120 849.150 78.540 ;
        RECT 858.185 78.355 921.630 78.975 ;
        RECT 922.640 77.910 979.410 78.405 ;
        RECT 981.610 78.120 1045.490 78.540 ;
        RECT 1054.525 78.355 1117.970 78.975 ;
        RECT 1118.965 77.915 1175.735 78.410 ;
        RECT 1177.950 78.120 1241.830 78.540 ;
        RECT 1250.865 78.355 1314.310 78.975 ;
        RECT 1.430 76.590 64.870 77.080 ;
        RECT 70.610 76.415 134.335 76.985 ;
        RECT 136.285 76.675 195.500 77.275 ;
        RECT 197.795 76.590 261.235 77.080 ;
        RECT 266.975 76.415 330.700 76.985 ;
        RECT 332.675 76.635 391.890 77.235 ;
        RECT 394.195 76.540 457.635 77.030 ;
        RECT 463.375 76.365 527.100 76.935 ;
        RECT 528.995 76.680 588.210 77.280 ;
        RECT 590.570 76.575 654.010 77.065 ;
        RECT 659.750 76.400 723.475 76.970 ;
        RECT 725.360 76.685 784.575 77.285 ;
        RECT 786.910 76.575 850.350 77.065 ;
        RECT 856.090 76.400 919.815 76.970 ;
        RECT 921.745 76.670 980.960 77.270 ;
        RECT 983.250 76.575 1046.690 77.065 ;
        RECT 1052.430 76.400 1116.155 76.970 ;
        RECT 1118.070 76.675 1177.285 77.275 ;
        RECT 1179.590 76.575 1243.030 77.065 ;
        RECT 1248.770 76.400 1312.495 76.970 ;
        RECT 1294.790 73.895 1310.810 74.305 ;
        RECT 101.380 73.325 103.975 73.755 ;
        RECT 297.745 73.325 300.340 73.755 ;
        RECT 494.145 73.275 496.740 73.705 ;
        RECT 690.520 73.310 693.115 73.740 ;
        RECT 886.860 73.310 889.455 73.740 ;
        RECT 1083.200 73.310 1085.795 73.740 ;
        RECT 1279.540 73.310 1282.135 73.740 ;
        RECT 1295.320 73.115 1310.800 73.570 ;
        RECT 102.060 72.200 119.430 72.540 ;
        RECT 298.425 72.200 315.795 72.540 ;
        RECT 494.825 72.150 512.195 72.490 ;
        RECT 691.200 72.185 708.570 72.525 ;
        RECT 887.540 72.185 904.910 72.525 ;
        RECT 1083.880 72.185 1101.250 72.525 ;
        RECT 1280.220 72.185 1297.590 72.525 ;
        RECT 34.130 70.420 36.835 70.760 ;
        RECT 230.495 70.420 233.200 70.760 ;
        RECT 426.895 70.370 429.600 70.710 ;
        RECT 623.270 70.405 625.975 70.745 ;
        RECT 819.610 70.405 822.315 70.745 ;
        RECT 1015.950 70.405 1018.655 70.745 ;
        RECT 1212.290 70.405 1214.995 70.745 ;
        RECT -0.280 69.175 5.700 69.320 ;
        RECT -4.160 69.015 5.700 69.175 ;
        RECT -4.160 68.880 0.070 69.015 ;
        RECT 18.395 69.005 21.140 69.335 ;
        RECT 195.925 69.185 202.065 69.320 ;
        RECT 192.010 69.015 202.065 69.185 ;
        RECT 192.010 68.890 196.240 69.015 ;
        RECT 214.760 69.005 217.505 69.335 ;
        RECT 588.635 69.305 588.950 69.325 ;
        RECT 392.315 69.270 392.630 69.280 ;
        RECT 392.315 69.145 398.465 69.270 ;
        RECT 388.400 68.965 398.465 69.145 ;
        RECT 388.400 68.850 392.630 68.965 ;
        RECT 411.160 68.955 413.905 69.285 ;
        RECT 588.635 69.190 594.840 69.305 ;
        RECT 584.720 69.000 594.840 69.190 ;
        RECT 584.720 68.895 588.950 69.000 ;
        RECT 607.535 68.990 610.280 69.320 ;
        RECT 785.000 69.305 785.315 69.330 ;
        RECT 785.000 69.195 791.180 69.305 ;
        RECT 781.085 69.000 791.180 69.195 ;
        RECT 781.085 68.900 785.315 69.000 ;
        RECT 803.875 68.990 806.620 69.320 ;
        RECT 981.385 69.305 981.700 69.315 ;
        RECT 981.385 69.180 987.520 69.305 ;
        RECT 977.470 69.000 987.520 69.180 ;
        RECT 977.470 68.885 981.700 69.000 ;
        RECT 1000.215 68.990 1002.960 69.320 ;
        RECT 1177.710 69.305 1178.025 69.320 ;
        RECT 1177.710 69.185 1183.860 69.305 ;
        RECT 1173.795 69.000 1183.860 69.185 ;
        RECT 1173.795 68.890 1178.025 69.000 ;
        RECT 1196.555 68.990 1199.300 69.320 ;
        RECT -0.265 68.500 5.680 68.575 ;
        RECT -2.265 68.280 5.680 68.500 ;
        RECT -2.265 68.155 0.050 68.280 ;
        RECT 18.400 68.255 21.140 68.585 ;
        RECT 196.015 68.510 202.045 68.575 ;
        RECT 193.905 68.280 202.045 68.510 ;
        RECT 193.905 68.165 196.220 68.280 ;
        RECT 214.765 68.255 217.505 68.585 ;
        RECT 392.285 68.470 398.445 68.525 ;
        RECT 390.295 68.230 398.445 68.470 ;
        RECT 390.295 68.125 392.610 68.230 ;
        RECT 411.165 68.205 413.905 68.535 ;
        RECT 588.620 68.515 594.820 68.560 ;
        RECT 586.615 68.265 594.820 68.515 ;
        RECT 586.615 68.170 588.930 68.265 ;
        RECT 607.540 68.240 610.280 68.570 ;
        RECT 784.985 68.560 785.295 68.565 ;
        RECT 784.985 68.520 791.160 68.560 ;
        RECT 782.980 68.265 791.160 68.520 ;
        RECT 782.980 68.175 785.295 68.265 ;
        RECT 803.880 68.240 806.620 68.570 ;
        RECT 981.555 68.550 987.500 68.560 ;
        RECT 981.370 68.505 987.500 68.550 ;
        RECT 979.365 68.265 987.500 68.505 ;
        RECT 979.365 68.160 981.680 68.265 ;
        RECT 1000.220 68.240 1002.960 68.570 ;
        RECT 1177.895 68.555 1183.840 68.560 ;
        RECT 1177.695 68.510 1183.840 68.555 ;
        RECT 1175.690 68.265 1183.840 68.510 ;
        RECT 1175.690 68.165 1178.005 68.265 ;
        RECT 1196.560 68.240 1199.300 68.570 ;
        RECT 1279.490 68.250 1281.515 68.635 ;
        RECT -3.420 67.855 5.715 67.860 ;
        RECT -3.745 67.725 5.715 67.855 ;
        RECT -55.980 67.565 5.715 67.725 ;
        RECT -55.980 67.555 -1.940 67.565 ;
        RECT -55.980 67.430 -3.520 67.555 ;
        RECT 18.405 67.235 36.130 67.555 ;
        RECT 116.585 67.230 119.430 67.610 ;
        RECT 192.945 67.565 202.080 67.860 ;
        RECT 214.770 67.235 232.495 67.555 ;
        RECT 312.950 67.230 315.795 67.610 ;
        RECT 389.345 67.515 398.480 67.810 ;
        RECT -3.300 67.095 5.670 67.230 ;
        RECT -55.235 66.935 5.670 67.095 ;
        RECT 193.065 66.935 202.035 67.230 ;
        RECT 411.170 67.185 428.895 67.505 ;
        RECT 509.350 67.180 512.195 67.560 ;
        RECT 585.720 67.550 594.855 67.845 ;
        RECT 607.545 67.220 625.270 67.540 ;
        RECT 705.725 67.215 708.570 67.595 ;
        RECT 782.060 67.550 791.195 67.845 ;
        RECT 803.885 67.220 821.610 67.540 ;
        RECT 902.065 67.215 904.910 67.595 ;
        RECT 978.400 67.550 987.535 67.845 ;
        RECT 1000.225 67.220 1017.950 67.540 ;
        RECT 1098.405 67.215 1101.250 67.595 ;
        RECT 1174.740 67.550 1183.875 67.845 ;
        RECT 1196.565 67.220 1214.290 67.540 ;
        RECT 1294.745 67.215 1297.590 67.595 ;
        RECT -55.235 66.790 -0.065 66.935 ;
        RECT 389.465 66.885 398.435 67.180 ;
        RECT 585.840 66.920 594.810 67.215 ;
        RECT 782.180 66.920 791.150 67.215 ;
        RECT 978.520 66.920 987.490 67.215 ;
        RECT 1174.860 66.920 1183.830 67.215 ;
        RECT -0.260 65.860 20.625 66.155 ;
        RECT 196.105 65.860 216.990 66.155 ;
        RECT 392.505 65.810 413.390 66.105 ;
        RECT 588.880 65.845 609.765 66.140 ;
        RECT 785.220 65.845 806.105 66.140 ;
        RECT 981.560 65.845 1002.445 66.140 ;
        RECT 1177.900 65.845 1198.785 66.140 ;
        RECT -0.260 64.995 21.210 65.290 ;
        RECT 33.820 65.115 37.720 65.600 ;
        RECT 116.560 65.155 118.845 65.580 ;
        RECT 196.105 64.995 217.575 65.290 ;
        RECT 230.185 65.115 234.085 65.600 ;
        RECT 312.925 65.155 315.210 65.580 ;
        RECT 392.505 64.945 413.975 65.240 ;
        RECT 426.585 65.065 430.485 65.550 ;
        RECT 509.325 65.105 511.610 65.530 ;
        RECT 588.880 64.980 610.350 65.275 ;
        RECT 622.960 65.100 626.860 65.585 ;
        RECT 705.700 65.140 707.985 65.565 ;
        RECT 785.220 64.980 806.690 65.275 ;
        RECT 819.300 65.100 823.200 65.585 ;
        RECT 902.040 65.140 904.325 65.565 ;
        RECT 981.560 64.980 1003.030 65.275 ;
        RECT 1015.640 65.100 1019.540 65.585 ;
        RECT 1098.380 65.140 1100.665 65.565 ;
        RECT 1177.900 64.980 1199.370 65.275 ;
        RECT 1211.980 65.100 1215.880 65.585 ;
        RECT 1279.655 65.300 1282.135 65.700 ;
        RECT 1294.720 65.140 1297.005 65.565 ;
        RECT 18.570 62.460 36.870 62.845 ;
        RECT 102.315 62.000 119.500 62.485 ;
        RECT 214.935 62.460 233.235 62.845 ;
        RECT 298.680 62.000 315.865 62.485 ;
        RECT 411.335 62.410 429.635 62.795 ;
        RECT 607.710 62.445 626.010 62.830 ;
        RECT 495.080 61.950 512.265 62.435 ;
        RECT 691.455 61.985 708.640 62.470 ;
        RECT 804.050 62.445 822.350 62.830 ;
        RECT 887.795 61.985 904.980 62.470 ;
        RECT 1000.390 62.445 1018.690 62.830 ;
        RECT 1084.135 61.985 1101.320 62.470 ;
        RECT 1196.730 62.445 1215.030 62.830 ;
        RECT 1280.475 61.985 1297.660 62.470 ;
        RECT 34.450 61.140 37.515 61.465 ;
        RECT 101.125 61.085 103.720 61.535 ;
        RECT 230.815 61.140 233.880 61.465 ;
        RECT 297.490 61.085 300.085 61.535 ;
        RECT 427.215 61.090 430.280 61.415 ;
        RECT 493.890 61.035 496.485 61.485 ;
        RECT 623.590 61.125 626.655 61.450 ;
        RECT 690.265 61.070 692.860 61.520 ;
        RECT 819.930 61.125 822.995 61.450 ;
        RECT 886.605 61.070 889.200 61.520 ;
        RECT 1016.270 61.125 1019.335 61.450 ;
        RECT 1082.945 61.070 1085.540 61.520 ;
        RECT 1212.610 61.125 1215.675 61.450 ;
        RECT 1279.285 61.070 1281.880 61.520 ;
        RECT -0.115 58.360 63.765 58.780 ;
        RECT 72.965 58.215 136.410 58.835 ;
        RECT 137.185 57.870 193.955 58.365 ;
        RECT 196.250 58.360 260.130 58.780 ;
        RECT 269.330 58.215 332.775 58.835 ;
        RECT 333.575 57.830 390.345 58.325 ;
        RECT 392.650 58.310 456.530 58.730 ;
        RECT 465.730 58.165 529.175 58.785 ;
        RECT 529.895 57.875 586.665 58.370 ;
        RECT 589.025 58.345 652.905 58.765 ;
        RECT 662.105 58.200 725.550 58.820 ;
        RECT 726.260 57.880 783.030 58.375 ;
        RECT 785.365 58.345 849.245 58.765 ;
        RECT 858.445 58.200 921.890 58.820 ;
        RECT 922.645 57.865 979.415 58.360 ;
        RECT 981.705 58.345 1045.585 58.765 ;
        RECT 1054.785 58.200 1118.230 58.820 ;
        RECT 1118.970 57.870 1175.740 58.365 ;
        RECT 1178.045 58.345 1241.925 58.765 ;
        RECT 1251.125 58.200 1314.570 58.820 ;
        RECT 1.525 56.815 64.965 57.305 ;
        RECT 70.870 56.260 134.595 56.830 ;
        RECT 136.290 56.630 195.505 57.230 ;
        RECT 197.890 56.815 261.330 57.305 ;
        RECT 267.235 56.260 330.960 56.830 ;
        RECT 332.680 56.590 391.895 57.190 ;
        RECT 394.290 56.765 457.730 57.255 ;
        RECT 463.635 56.210 527.360 56.780 ;
        RECT 529.000 56.635 588.215 57.235 ;
        RECT 590.665 56.800 654.105 57.290 ;
        RECT 660.010 56.245 723.735 56.815 ;
        RECT 725.365 56.640 784.580 57.240 ;
        RECT 787.005 56.800 850.445 57.290 ;
        RECT 856.350 56.245 920.075 56.815 ;
        RECT 921.750 56.625 980.965 57.225 ;
        RECT 983.345 56.800 1046.785 57.290 ;
        RECT 1052.690 56.245 1116.415 56.815 ;
        RECT 1118.075 56.630 1177.290 57.230 ;
        RECT 1179.685 56.800 1243.125 57.290 ;
        RECT 1249.030 56.245 1312.755 56.815 ;
        RECT 1294.790 53.925 1310.810 54.335 ;
        RECT 101.380 53.355 103.975 53.785 ;
        RECT 297.745 53.355 300.340 53.785 ;
        RECT 494.145 53.305 496.740 53.735 ;
        RECT 690.520 53.340 693.115 53.770 ;
        RECT 886.860 53.340 889.455 53.770 ;
        RECT 1083.200 53.340 1085.795 53.770 ;
        RECT 1279.540 53.340 1282.135 53.770 ;
        RECT 1295.320 53.145 1310.800 53.600 ;
        RECT 102.060 52.230 119.430 52.570 ;
        RECT 298.425 52.230 315.795 52.570 ;
        RECT 494.825 52.180 512.195 52.520 ;
        RECT 691.200 52.215 708.570 52.555 ;
        RECT 887.540 52.215 904.910 52.555 ;
        RECT 1083.880 52.215 1101.250 52.555 ;
        RECT 1280.220 52.215 1297.590 52.555 ;
        RECT 34.080 50.610 36.785 50.950 ;
        RECT 230.445 50.610 233.150 50.950 ;
        RECT 426.845 50.560 429.550 50.900 ;
        RECT 623.220 50.595 625.925 50.935 ;
        RECT 819.560 50.595 822.265 50.935 ;
        RECT 1015.900 50.595 1018.605 50.935 ;
        RECT 1212.240 50.595 1214.945 50.935 ;
        RECT -0.330 49.455 5.650 49.510 ;
        RECT -4.090 49.205 5.650 49.455 ;
        RECT -4.090 49.160 0.140 49.205 ;
        RECT 18.345 49.195 21.090 49.525 ;
        RECT 196.035 49.465 202.015 49.510 ;
        RECT 192.080 49.205 202.015 49.465 ;
        RECT 192.080 49.170 196.310 49.205 ;
        RECT 214.710 49.195 217.455 49.525 ;
        RECT 392.435 49.425 398.415 49.460 ;
        RECT 388.470 49.155 398.415 49.425 ;
        RECT 388.470 49.130 392.700 49.155 ;
        RECT 411.110 49.145 413.855 49.475 ;
        RECT 588.810 49.470 594.790 49.495 ;
        RECT 584.790 49.190 594.790 49.470 ;
        RECT 584.790 49.175 589.020 49.190 ;
        RECT 607.485 49.180 610.230 49.510 ;
        RECT 785.150 49.475 791.130 49.495 ;
        RECT 781.155 49.190 791.130 49.475 ;
        RECT 781.155 49.180 785.385 49.190 ;
        RECT 803.825 49.180 806.570 49.510 ;
        RECT 981.490 49.460 987.470 49.495 ;
        RECT 977.540 49.190 987.470 49.460 ;
        RECT 977.540 49.165 981.770 49.190 ;
        RECT 1000.165 49.180 1002.910 49.510 ;
        RECT 1177.830 49.465 1183.810 49.495 ;
        RECT 1173.865 49.190 1183.810 49.465 ;
        RECT 1173.865 49.170 1178.095 49.190 ;
        RECT 1196.505 49.180 1199.250 49.510 ;
        RECT -2.195 48.765 0.120 48.780 ;
        RECT -2.195 48.470 5.630 48.765 ;
        RECT -2.195 48.435 0.120 48.470 ;
        RECT 18.350 48.445 21.090 48.775 ;
        RECT 193.975 48.765 196.290 48.790 ;
        RECT 193.975 48.470 201.995 48.765 ;
        RECT 193.975 48.445 196.290 48.470 ;
        RECT 214.715 48.445 217.455 48.775 ;
        RECT 586.685 48.750 589.000 48.795 ;
        RECT 390.365 48.715 392.680 48.750 ;
        RECT 390.365 48.420 398.395 48.715 ;
        RECT 390.365 48.405 392.680 48.420 ;
        RECT 411.115 48.395 413.855 48.725 ;
        RECT 586.685 48.455 594.770 48.750 ;
        RECT 586.685 48.450 589.000 48.455 ;
        RECT 607.490 48.430 610.230 48.760 ;
        RECT 783.050 48.750 785.365 48.800 ;
        RECT 783.050 48.455 791.110 48.750 ;
        RECT 803.830 48.430 806.570 48.760 ;
        RECT 979.435 48.750 981.750 48.785 ;
        RECT 979.435 48.455 987.450 48.750 ;
        RECT 979.435 48.440 981.750 48.455 ;
        RECT 1000.170 48.430 1002.910 48.760 ;
        RECT 1175.760 48.750 1178.075 48.790 ;
        RECT 1175.760 48.455 1183.790 48.750 ;
        RECT 1175.760 48.445 1178.075 48.455 ;
        RECT 1196.510 48.430 1199.250 48.760 ;
        RECT 1279.490 48.280 1281.515 48.665 ;
        RECT -3.470 48.005 5.665 48.050 ;
        RECT -55.895 47.755 5.665 48.005 ;
        RECT 192.895 47.755 202.030 48.050 ;
        RECT -55.895 47.710 0.055 47.755 ;
        RECT 18.355 47.425 36.080 47.745 ;
        RECT -3.350 47.375 5.620 47.420 ;
        RECT -55.140 47.125 5.620 47.375 ;
        RECT 116.585 47.260 119.430 47.640 ;
        RECT 214.720 47.425 232.445 47.745 ;
        RECT 389.295 47.705 398.430 48.000 ;
        RECT 585.670 47.740 594.805 48.035 ;
        RECT 782.010 47.740 791.145 48.035 ;
        RECT 978.350 47.740 987.485 48.035 ;
        RECT 1174.690 47.740 1183.825 48.035 ;
        RECT 193.015 47.125 201.985 47.420 ;
        RECT 312.950 47.260 315.795 47.640 ;
        RECT 411.120 47.375 428.845 47.695 ;
        RECT -55.140 47.070 0.005 47.125 ;
        RECT 389.415 47.075 398.385 47.370 ;
        RECT 509.350 47.210 512.195 47.590 ;
        RECT 607.495 47.410 625.220 47.730 ;
        RECT 585.790 47.110 594.760 47.405 ;
        RECT 705.725 47.245 708.570 47.625 ;
        RECT 803.835 47.410 821.560 47.730 ;
        RECT 782.130 47.110 791.100 47.405 ;
        RECT 902.065 47.245 904.910 47.625 ;
        RECT 1000.175 47.410 1017.900 47.730 ;
        RECT 978.470 47.110 987.440 47.405 ;
        RECT 1098.405 47.245 1101.250 47.625 ;
        RECT 1196.515 47.410 1214.240 47.730 ;
        RECT 1174.810 47.110 1183.780 47.405 ;
        RECT 1294.745 47.245 1297.590 47.625 ;
        RECT -0.310 46.050 20.575 46.345 ;
        RECT 196.055 46.050 216.940 46.345 ;
        RECT 392.455 46.000 413.340 46.295 ;
        RECT 588.830 46.035 609.715 46.330 ;
        RECT 785.170 46.035 806.055 46.330 ;
        RECT 981.510 46.035 1002.395 46.330 ;
        RECT 1177.850 46.035 1198.735 46.330 ;
        RECT -0.310 45.185 21.160 45.480 ;
        RECT 33.770 45.305 37.670 45.790 ;
        RECT 116.560 45.185 118.845 45.610 ;
        RECT 196.055 45.185 217.525 45.480 ;
        RECT 230.135 45.305 234.035 45.790 ;
        RECT 312.925 45.185 315.210 45.610 ;
        RECT 392.455 45.135 413.925 45.430 ;
        RECT 426.535 45.255 430.435 45.740 ;
        RECT 509.325 45.135 511.610 45.560 ;
        RECT 588.830 45.170 610.300 45.465 ;
        RECT 622.910 45.290 626.810 45.775 ;
        RECT 705.700 45.170 707.985 45.595 ;
        RECT 785.170 45.170 806.640 45.465 ;
        RECT 819.250 45.290 823.150 45.775 ;
        RECT 902.040 45.170 904.325 45.595 ;
        RECT 981.510 45.170 1002.980 45.465 ;
        RECT 1015.590 45.290 1019.490 45.775 ;
        RECT 1098.380 45.170 1100.665 45.595 ;
        RECT 1177.850 45.170 1199.320 45.465 ;
        RECT 1211.930 45.290 1215.830 45.775 ;
        RECT 1279.655 45.330 1282.135 45.730 ;
        RECT 1294.720 45.170 1297.005 45.595 ;
        RECT 18.520 42.650 36.820 43.035 ;
        RECT 214.885 42.650 233.185 43.035 ;
        RECT 411.285 42.600 429.585 42.985 ;
        RECT 607.660 42.635 625.960 43.020 ;
        RECT 804.000 42.635 822.300 43.020 ;
        RECT 1000.340 42.635 1018.640 43.020 ;
        RECT 1196.680 42.635 1214.980 43.020 ;
        RECT 102.315 42.030 119.500 42.515 ;
        RECT 298.680 42.030 315.865 42.515 ;
        RECT 495.080 41.980 512.265 42.465 ;
        RECT 691.455 42.015 708.640 42.500 ;
        RECT 887.795 42.015 904.980 42.500 ;
        RECT 1084.135 42.015 1101.320 42.500 ;
        RECT 1280.475 42.015 1297.660 42.500 ;
        RECT 34.400 41.330 37.465 41.655 ;
        RECT 101.125 41.115 103.720 41.565 ;
        RECT 230.765 41.330 233.830 41.655 ;
        RECT 297.490 41.115 300.085 41.565 ;
        RECT 427.165 41.280 430.230 41.605 ;
        RECT 493.890 41.065 496.485 41.515 ;
        RECT 623.540 41.315 626.605 41.640 ;
        RECT 690.265 41.100 692.860 41.550 ;
        RECT 819.880 41.315 822.945 41.640 ;
        RECT 886.605 41.100 889.200 41.550 ;
        RECT 1016.220 41.315 1019.285 41.640 ;
        RECT 1082.945 41.100 1085.540 41.550 ;
        RECT 1212.560 41.315 1215.625 41.640 ;
        RECT 1279.285 41.100 1281.880 41.550 ;
        RECT -0.115 38.550 63.765 38.970 ;
        RECT 73.075 38.325 136.520 38.945 ;
        RECT 137.190 38.205 193.960 38.700 ;
        RECT 196.250 38.550 260.130 38.970 ;
        RECT 269.440 38.325 332.885 38.945 ;
        RECT 333.580 38.165 390.350 38.660 ;
        RECT 392.650 38.500 456.530 38.920 ;
        RECT 465.840 38.275 529.285 38.895 ;
        RECT 529.900 38.210 586.670 38.705 ;
        RECT 589.025 38.535 652.905 38.955 ;
        RECT 662.215 38.310 725.660 38.930 ;
        RECT 726.265 38.215 783.035 38.710 ;
        RECT 785.365 38.535 849.245 38.955 ;
        RECT 858.555 38.310 922.000 38.930 ;
        RECT 922.650 38.200 979.420 38.695 ;
        RECT 981.705 38.535 1045.585 38.955 ;
        RECT 1054.895 38.310 1118.340 38.930 ;
        RECT 1118.975 38.205 1175.745 38.700 ;
        RECT 1178.045 38.535 1241.925 38.955 ;
        RECT 1251.235 38.310 1314.680 38.930 ;
        RECT 1.525 37.005 64.965 37.495 ;
        RECT 136.295 36.965 195.510 37.565 ;
        RECT 197.890 37.005 261.330 37.495 ;
        RECT 70.980 36.370 134.705 36.940 ;
        RECT 267.345 36.370 331.070 36.940 ;
        RECT 332.685 36.925 391.900 37.525 ;
        RECT 394.290 36.955 457.730 37.445 ;
        RECT 529.005 36.970 588.220 37.570 ;
        RECT 590.665 36.990 654.105 37.480 ;
        RECT 725.370 36.975 784.585 37.575 ;
        RECT 787.005 36.990 850.445 37.480 ;
        RECT 921.755 36.960 980.970 37.560 ;
        RECT 983.345 36.990 1046.785 37.480 ;
        RECT 1118.080 36.965 1177.295 37.565 ;
        RECT 1179.685 36.990 1243.125 37.480 ;
        RECT 463.745 36.320 527.470 36.890 ;
        RECT 660.120 36.355 723.845 36.925 ;
        RECT 856.460 36.355 920.185 36.925 ;
        RECT 1052.800 36.355 1116.525 36.925 ;
        RECT 1249.140 36.355 1312.865 36.925 ;
        RECT 1294.790 34.260 1310.810 34.670 ;
        RECT 101.380 33.690 103.975 34.120 ;
        RECT 297.745 33.690 300.340 34.120 ;
        RECT 494.145 33.640 496.740 34.070 ;
        RECT 690.520 33.675 693.115 34.105 ;
        RECT 886.860 33.675 889.455 34.105 ;
        RECT 1083.200 33.675 1085.795 34.105 ;
        RECT 1279.540 33.675 1282.135 34.105 ;
        RECT 1295.320 33.480 1310.800 33.935 ;
        RECT 102.060 32.565 119.430 32.905 ;
        RECT 298.425 32.565 315.795 32.905 ;
        RECT 494.825 32.515 512.195 32.855 ;
        RECT 691.200 32.550 708.570 32.890 ;
        RECT 887.540 32.550 904.910 32.890 ;
        RECT 1083.880 32.550 1101.250 32.890 ;
        RECT 1280.220 32.550 1297.590 32.890 ;
        RECT 230.415 30.815 233.120 31.155 ;
        RECT 426.815 30.765 429.520 31.105 ;
        RECT 623.190 30.800 625.895 31.140 ;
        RECT 819.530 30.800 822.235 31.140 ;
        RECT 1015.870 30.800 1018.575 31.140 ;
        RECT 1212.210 30.800 1214.915 31.140 ;
        RECT 196.005 29.655 201.985 29.715 ;
        RECT 192.085 29.410 201.985 29.655 ;
        RECT 192.085 29.360 196.315 29.410 ;
        RECT 214.680 29.400 217.425 29.730 ;
        RECT 392.405 29.615 398.385 29.665 ;
        RECT 388.475 29.360 398.385 29.615 ;
        RECT 388.475 29.320 392.705 29.360 ;
        RECT 411.080 29.350 413.825 29.680 ;
        RECT 588.780 29.660 594.760 29.700 ;
        RECT 584.795 29.395 594.760 29.660 ;
        RECT 584.795 29.365 589.025 29.395 ;
        RECT 607.455 29.385 610.200 29.715 ;
        RECT 785.120 29.665 791.100 29.700 ;
        RECT 781.160 29.395 791.100 29.665 ;
        RECT 781.160 29.370 785.390 29.395 ;
        RECT 803.795 29.385 806.540 29.715 ;
        RECT 981.460 29.650 987.440 29.700 ;
        RECT 977.545 29.395 987.440 29.650 ;
        RECT 977.545 29.355 981.775 29.395 ;
        RECT 1000.135 29.385 1002.880 29.715 ;
        RECT 1177.800 29.655 1183.780 29.700 ;
        RECT 1173.870 29.395 1183.780 29.655 ;
        RECT 1173.870 29.360 1178.100 29.395 ;
        RECT 1196.475 29.385 1199.220 29.715 ;
        RECT 193.980 28.970 196.295 28.980 ;
        RECT 193.980 28.675 201.965 28.970 ;
        RECT 193.980 28.635 196.295 28.675 ;
        RECT 214.685 28.650 217.425 28.980 ;
        RECT 586.690 28.955 589.005 28.985 ;
        RECT 390.370 28.920 392.685 28.940 ;
        RECT 390.370 28.625 398.365 28.920 ;
        RECT 390.370 28.595 392.685 28.625 ;
        RECT 411.085 28.600 413.825 28.930 ;
        RECT 586.690 28.660 594.740 28.955 ;
        RECT 586.690 28.640 589.005 28.660 ;
        RECT 607.460 28.635 610.200 28.965 ;
        RECT 783.055 28.955 785.370 28.990 ;
        RECT 783.055 28.660 791.080 28.955 ;
        RECT 783.055 28.645 785.370 28.660 ;
        RECT 803.800 28.635 806.540 28.965 ;
        RECT 979.440 28.955 981.755 28.975 ;
        RECT 979.440 28.660 987.420 28.955 ;
        RECT 979.440 28.630 981.755 28.660 ;
        RECT 1000.140 28.635 1002.880 28.965 ;
        RECT 1175.765 28.955 1178.080 28.980 ;
        RECT 1175.765 28.660 1183.760 28.955 ;
        RECT 1175.765 28.635 1178.080 28.660 ;
        RECT 1196.480 28.635 1199.220 28.965 ;
        RECT 1279.490 28.615 1281.515 29.000 ;
        RECT -3.500 28.250 5.635 28.255 ;
        RECT -3.620 28.195 5.635 28.250 ;
        RECT -55.875 27.960 5.635 28.195 ;
        RECT -55.875 27.900 -3.460 27.960 ;
        RECT 18.325 27.630 36.050 27.950 ;
        RECT -3.380 27.565 5.590 27.625 ;
        RECT 116.585 27.595 119.430 27.975 ;
        RECT 192.865 27.960 202.000 28.255 ;
        RECT 214.690 27.630 232.415 27.950 ;
        RECT -55.130 27.330 5.590 27.565 ;
        RECT 192.985 27.330 201.955 27.625 ;
        RECT 312.950 27.595 315.795 27.975 ;
        RECT 389.265 27.910 398.400 28.205 ;
        RECT 585.640 27.945 594.775 28.240 ;
        RECT 411.090 27.580 428.815 27.900 ;
        RECT -55.130 27.260 0.010 27.330 ;
        RECT 389.385 27.280 398.355 27.575 ;
        RECT 509.350 27.545 512.195 27.925 ;
        RECT 607.465 27.615 625.190 27.935 ;
        RECT 585.760 27.315 594.730 27.610 ;
        RECT 705.725 27.580 708.570 27.960 ;
        RECT 781.980 27.945 791.115 28.240 ;
        RECT 803.805 27.615 821.530 27.935 ;
        RECT 782.100 27.315 791.070 27.610 ;
        RECT 902.065 27.580 904.910 27.960 ;
        RECT 978.320 27.945 987.455 28.240 ;
        RECT 1000.145 27.615 1017.870 27.935 ;
        RECT 978.440 27.315 987.410 27.610 ;
        RECT 1098.405 27.580 1101.250 27.960 ;
        RECT 1174.660 27.945 1183.795 28.240 ;
        RECT 1196.485 27.615 1214.210 27.935 ;
        RECT 1174.780 27.315 1183.750 27.610 ;
        RECT 1294.745 27.580 1297.590 27.960 ;
        RECT -0.340 26.255 20.545 26.550 ;
        RECT 196.025 26.255 216.910 26.550 ;
        RECT 392.425 26.205 413.310 26.500 ;
        RECT 588.800 26.240 609.685 26.535 ;
        RECT 785.140 26.240 806.025 26.535 ;
        RECT 981.480 26.240 1002.365 26.535 ;
        RECT 1177.820 26.240 1198.705 26.535 ;
        RECT -0.340 25.390 21.130 25.685 ;
        RECT 33.740 25.510 37.640 25.995 ;
        RECT 116.560 25.520 118.845 25.945 ;
        RECT 196.025 25.390 217.495 25.685 ;
        RECT 230.105 25.510 234.005 25.995 ;
        RECT 312.925 25.520 315.210 25.945 ;
        RECT 392.425 25.340 413.895 25.635 ;
        RECT 426.505 25.460 430.405 25.945 ;
        RECT 509.325 25.470 511.610 25.895 ;
        RECT 588.800 25.375 610.270 25.670 ;
        RECT 622.880 25.495 626.780 25.980 ;
        RECT 705.700 25.505 707.985 25.930 ;
        RECT 785.140 25.375 806.610 25.670 ;
        RECT 819.220 25.495 823.120 25.980 ;
        RECT 902.040 25.505 904.325 25.930 ;
        RECT 981.480 25.375 1002.950 25.670 ;
        RECT 1015.560 25.495 1019.460 25.980 ;
        RECT 1098.380 25.505 1100.665 25.930 ;
        RECT 1177.820 25.375 1199.290 25.670 ;
        RECT 1211.900 25.495 1215.800 25.980 ;
        RECT 1279.655 25.665 1282.135 26.065 ;
        RECT 1294.720 25.505 1297.005 25.930 ;
        RECT 18.490 22.855 36.790 23.240 ;
        RECT 214.855 22.855 233.155 23.240 ;
        RECT 102.315 22.365 119.500 22.850 ;
        RECT 298.680 22.365 315.865 22.850 ;
        RECT 411.255 22.805 429.555 23.190 ;
        RECT 607.630 22.840 625.930 23.225 ;
        RECT 803.970 22.840 822.270 23.225 ;
        RECT 1000.310 22.840 1018.610 23.225 ;
        RECT 1196.650 22.840 1214.950 23.225 ;
        RECT 495.080 22.315 512.265 22.800 ;
        RECT 691.455 22.350 708.640 22.835 ;
        RECT 887.795 22.350 904.980 22.835 ;
        RECT 1084.135 22.350 1101.320 22.835 ;
        RECT 1280.475 22.350 1297.660 22.835 ;
        RECT 34.370 21.535 37.435 21.860 ;
        RECT 101.125 21.450 103.720 21.900 ;
        RECT 230.735 21.535 233.800 21.860 ;
        RECT 297.490 21.450 300.085 21.900 ;
        RECT 427.135 21.485 430.200 21.810 ;
        RECT 493.890 21.400 496.485 21.850 ;
        RECT 623.510 21.520 626.575 21.845 ;
        RECT 690.265 21.435 692.860 21.885 ;
        RECT 819.850 21.520 822.915 21.845 ;
        RECT 886.605 21.435 889.200 21.885 ;
        RECT 1016.190 21.520 1019.255 21.845 ;
        RECT 1082.945 21.435 1085.540 21.885 ;
        RECT 1212.530 21.520 1215.595 21.845 ;
        RECT 1279.285 21.435 1281.880 21.885 ;
        RECT 87.895 7.890 195.410 8.185 ;
        RECT 284.290 7.900 391.805 8.195 ;
        RECT 480.610 7.845 588.125 8.140 ;
        RECT 676.975 7.885 784.490 8.180 ;
        RECT 873.360 7.885 980.875 8.180 ;
        RECT 1069.685 7.890 1177.200 8.185 ;
        RECT 87.905 5.825 194.190 6.170 ;
        RECT 284.300 5.825 390.585 6.170 ;
        RECT 480.650 5.775 586.935 6.120 ;
        RECT 677.020 5.810 783.305 6.155 ;
        RECT 873.405 5.795 979.690 6.140 ;
        RECT 1069.730 5.800 1176.015 6.145 ;
  END
END 8b_mult
END LIBRARY

