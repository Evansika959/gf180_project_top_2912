VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fa16b_rev
  CLASS BLOCK ;
  FOREIGN fa16b_rev ;
  ORIGIN -80.625 184.225 ;
  SIZE 1.120 BY 15.925 ;
  PIN s15
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 115.190 -153.920 115.570 -153.540 ;
        RECT 112.515 -154.345 114.255 -154.055 ;
        RECT 113.870 -158.940 124.275 -158.605 ;
        RECT 113.840 -160.260 115.620 -159.970 ;
        RECT 112.570 -160.875 112.950 -160.495 ;
      LAYER Metal2 ;
        RECT 112.600 -160.935 112.900 -154.005 ;
        RECT 113.910 -160.335 114.210 -153.985 ;
        RECT 115.225 -160.305 115.520 -153.480 ;
    END
  END s15
  PIN s15_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 122.090 -153.930 122.470 -153.550 ;
        RECT 119.015 -154.425 121.640 -154.015 ;
        RECT 121.200 -156.865 124.275 -156.590 ;
        RECT 121.215 -160.290 122.525 -159.970 ;
        RECT 119.025 -160.845 119.405 -160.465 ;
      LAYER Metal2 ;
        RECT 119.065 -160.935 119.365 -153.995 ;
        RECT 121.275 -160.360 121.555 -154.000 ;
        RECT 122.125 -160.360 122.425 -153.540 ;
    END
  END s15_not
  PIN s14
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 115.190 -134.255 115.570 -133.875 ;
        RECT 112.515 -134.680 114.255 -134.390 ;
        RECT 113.870 -139.275 124.275 -138.940 ;
        RECT 113.840 -140.595 115.620 -140.305 ;
        RECT 112.570 -141.210 112.950 -140.830 ;
      LAYER Metal2 ;
        RECT 112.600 -141.270 112.900 -134.340 ;
        RECT 113.910 -140.670 114.210 -134.320 ;
        RECT 115.225 -140.640 115.520 -133.815 ;
    END
  END s14
  PIN s14_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 122.090 -134.265 122.470 -133.885 ;
        RECT 119.015 -134.760 121.640 -134.350 ;
        RECT 121.200 -137.200 124.275 -136.925 ;
        RECT 121.215 -140.625 122.525 -140.305 ;
        RECT 119.025 -141.180 119.405 -140.800 ;
      LAYER Metal2 ;
        RECT 119.065 -141.270 119.365 -134.330 ;
        RECT 121.275 -140.695 121.555 -134.335 ;
        RECT 122.125 -140.695 122.425 -133.875 ;
    END
  END s14_not
  PIN s13
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 115.190 -114.285 115.570 -113.905 ;
        RECT 112.515 -114.710 114.255 -114.420 ;
        RECT 113.870 -119.305 124.275 -118.970 ;
        RECT 113.840 -120.625 115.620 -120.335 ;
        RECT 112.570 -121.240 112.950 -120.860 ;
      LAYER Metal2 ;
        RECT 112.600 -121.300 112.900 -114.370 ;
        RECT 113.910 -120.700 114.210 -114.350 ;
        RECT 115.225 -120.670 115.520 -113.845 ;
    END
  END s13
  PIN s13_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 122.090 -114.295 122.470 -113.915 ;
        RECT 119.015 -114.790 121.640 -114.380 ;
        RECT 121.200 -117.230 124.275 -116.955 ;
        RECT 121.215 -120.655 122.525 -120.335 ;
        RECT 119.025 -121.210 119.405 -120.830 ;
      LAYER Metal2 ;
        RECT 119.065 -121.300 119.365 -114.360 ;
        RECT 121.275 -120.725 121.555 -114.365 ;
        RECT 122.125 -120.725 122.425 -113.905 ;
    END
  END s13_not
  PIN s12
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 115.085 -94.570 115.465 -94.190 ;
        RECT 112.410 -94.995 114.150 -94.705 ;
        RECT 113.765 -99.590 124.170 -99.255 ;
        RECT 113.735 -100.910 115.515 -100.620 ;
        RECT 112.465 -101.525 112.845 -101.145 ;
      LAYER Metal2 ;
        RECT 112.495 -101.585 112.795 -94.655 ;
        RECT 113.805 -100.985 114.105 -94.635 ;
        RECT 115.120 -100.955 115.415 -94.130 ;
    END
  END s12
  PIN s12_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 121.985 -94.580 122.365 -94.200 ;
        RECT 118.910 -95.075 121.535 -94.665 ;
        RECT 121.095 -97.515 124.170 -97.240 ;
        RECT 121.110 -100.940 122.420 -100.620 ;
        RECT 118.920 -101.495 119.300 -101.115 ;
      LAYER Metal2 ;
        RECT 118.960 -101.585 119.260 -94.645 ;
        RECT 121.170 -101.010 121.450 -94.650 ;
        RECT 122.020 -101.010 122.320 -94.190 ;
    END
  END s12_not
  PIN s11
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 115.165 -74.815 115.545 -74.435 ;
        RECT 112.490 -75.240 114.230 -74.950 ;
        RECT 113.845 -79.835 124.250 -79.500 ;
        RECT 113.815 -81.155 115.595 -80.865 ;
        RECT 112.545 -81.770 112.925 -81.390 ;
      LAYER Metal2 ;
        RECT 112.575 -81.830 112.875 -74.900 ;
        RECT 113.885 -81.230 114.185 -74.880 ;
        RECT 115.200 -81.200 115.495 -74.375 ;
    END
  END s11
  PIN s11_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 122.065 -74.825 122.445 -74.445 ;
        RECT 118.990 -75.320 121.615 -74.910 ;
        RECT 121.175 -77.760 124.250 -77.485 ;
        RECT 121.190 -81.185 122.500 -80.865 ;
        RECT 119.000 -81.740 119.380 -81.360 ;
      LAYER Metal2 ;
        RECT 119.040 -81.830 119.340 -74.890 ;
        RECT 121.250 -81.255 121.530 -74.895 ;
        RECT 122.100 -81.255 122.400 -74.435 ;
    END
  END s11_not
  PIN s10
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 115.165 -55.020 115.545 -54.640 ;
        RECT 112.490 -55.445 114.230 -55.155 ;
        RECT 113.845 -60.040 124.250 -59.705 ;
        RECT 113.815 -61.360 115.595 -61.070 ;
        RECT 112.545 -61.975 112.925 -61.595 ;
      LAYER Metal2 ;
        RECT 112.575 -62.035 112.875 -55.105 ;
        RECT 113.885 -61.435 114.185 -55.085 ;
        RECT 115.200 -61.405 115.495 -54.580 ;
    END
  END s10
  PIN s10_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 122.065 -55.030 122.445 -54.650 ;
        RECT 118.990 -55.525 121.615 -55.115 ;
        RECT 121.175 -57.965 124.250 -57.690 ;
        RECT 121.190 -61.390 122.500 -61.070 ;
        RECT 119.000 -61.945 119.380 -61.565 ;
      LAYER Metal2 ;
        RECT 119.040 -62.035 119.340 -55.095 ;
        RECT 121.250 -61.460 121.530 -55.100 ;
        RECT 122.100 -61.460 122.400 -54.640 ;
    END
  END s10_not
  PIN s4
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 115.065 63.540 115.445 63.920 ;
        RECT 112.390 63.115 114.130 63.405 ;
        RECT 113.745 58.520 124.150 58.855 ;
        RECT 113.715 57.200 115.495 57.490 ;
        RECT 112.445 56.585 112.825 56.965 ;
      LAYER Metal2 ;
        RECT 112.475 56.525 112.775 63.455 ;
        RECT 113.785 57.125 114.085 63.475 ;
        RECT 115.100 57.155 115.395 63.980 ;
    END
  END s4
  PIN s4_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 121.965 63.530 122.345 63.910 ;
        RECT 118.890 63.035 121.515 63.445 ;
        RECT 121.075 60.595 124.150 60.870 ;
        RECT 121.090 57.170 122.400 57.490 ;
        RECT 118.900 56.615 119.280 56.995 ;
      LAYER Metal2 ;
        RECT 118.940 56.525 119.240 63.465 ;
        RECT 121.150 57.100 121.430 63.460 ;
        RECT 122.000 57.100 122.300 63.920 ;
    END
  END s4_not
  PIN s9
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 115.010 -35.375 115.390 -34.995 ;
        RECT 112.335 -35.800 114.075 -35.510 ;
        RECT 113.690 -40.395 124.095 -40.060 ;
        RECT 113.660 -41.715 115.440 -41.425 ;
        RECT 112.390 -42.330 112.770 -41.950 ;
      LAYER Metal2 ;
        RECT 112.420 -42.390 112.720 -35.460 ;
        RECT 113.730 -41.790 114.030 -35.440 ;
        RECT 115.045 -41.760 115.340 -34.935 ;
    END
  END s9
  PIN s9_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 121.910 -35.385 122.290 -35.005 ;
        RECT 118.835 -35.880 121.460 -35.470 ;
        RECT 121.020 -38.320 124.095 -38.045 ;
        RECT 121.035 -41.745 122.345 -41.425 ;
        RECT 118.845 -42.300 119.225 -41.920 ;
      LAYER Metal2 ;
        RECT 118.885 -42.390 119.185 -35.450 ;
        RECT 121.095 -41.815 121.375 -35.455 ;
        RECT 121.945 -41.815 122.245 -34.995 ;
    END
  END s9_not
  PIN s3
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 115.145 83.295 115.525 83.675 ;
        RECT 112.470 82.870 114.210 83.160 ;
        RECT 113.825 78.275 124.230 78.610 ;
        RECT 113.795 76.955 115.575 77.245 ;
        RECT 112.525 76.340 112.905 76.720 ;
      LAYER Metal2 ;
        RECT 112.555 76.280 112.855 83.210 ;
        RECT 113.865 76.880 114.165 83.230 ;
        RECT 115.180 76.910 115.475 83.735 ;
    END
  END s3
  PIN s3_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 122.045 83.285 122.425 83.665 ;
        RECT 118.970 82.790 121.595 83.200 ;
        RECT 121.155 80.350 124.230 80.625 ;
        RECT 121.170 76.925 122.480 77.245 ;
        RECT 118.980 76.370 119.360 76.750 ;
      LAYER Metal2 ;
        RECT 119.020 76.280 119.320 83.220 ;
        RECT 121.230 76.855 121.510 83.215 ;
        RECT 122.080 76.855 122.380 83.675 ;
    END
  END s3_not
  PIN s8
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 115.210 -15.650 115.590 -15.270 ;
        RECT 112.535 -16.075 114.275 -15.785 ;
        RECT 113.890 -20.670 124.295 -20.335 ;
        RECT 113.860 -21.990 115.640 -21.700 ;
        RECT 112.590 -22.605 112.970 -22.225 ;
      LAYER Metal2 ;
        RECT 112.620 -22.665 112.920 -15.735 ;
        RECT 113.930 -22.065 114.230 -15.715 ;
        RECT 115.245 -22.035 115.540 -15.210 ;
    END
  END s8
  PIN s8_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 122.110 -15.660 122.490 -15.280 ;
        RECT 119.035 -16.155 121.660 -15.745 ;
        RECT 121.220 -18.595 124.295 -18.320 ;
        RECT 121.235 -22.020 122.545 -21.700 ;
        RECT 119.045 -22.575 119.425 -22.195 ;
      LAYER Metal2 ;
        RECT 119.085 -22.665 119.385 -15.725 ;
        RECT 121.295 -22.090 121.575 -15.730 ;
        RECT 122.145 -22.090 122.445 -15.270 ;
    END
  END s8_not
  PIN s2
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 115.145 103.090 115.525 103.470 ;
        RECT 112.470 102.665 114.210 102.955 ;
        RECT 113.825 98.070 124.230 98.405 ;
        RECT 113.795 96.750 115.575 97.040 ;
        RECT 112.525 96.135 112.905 96.515 ;
      LAYER Metal2 ;
        RECT 112.555 96.075 112.855 103.005 ;
        RECT 113.865 96.675 114.165 103.025 ;
        RECT 115.180 96.705 115.475 103.530 ;
    END
  END s2
  PIN s2_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 122.045 103.080 122.425 103.460 ;
        RECT 118.970 102.585 121.595 102.995 ;
        RECT 121.155 100.145 124.230 100.420 ;
        RECT 121.170 96.720 122.480 97.040 ;
        RECT 118.980 96.165 119.360 96.545 ;
      LAYER Metal2 ;
        RECT 119.020 96.075 119.320 103.015 ;
        RECT 121.230 96.650 121.510 103.010 ;
        RECT 122.080 96.650 122.380 103.470 ;
    END
  END s2_not
  PIN s7
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 115.170 4.190 115.550 4.570 ;
        RECT 112.495 3.765 114.235 4.055 ;
        RECT 113.850 -0.830 124.255 -0.495 ;
        RECT 113.820 -2.150 115.600 -1.860 ;
        RECT 112.550 -2.765 112.930 -2.385 ;
      LAYER Metal2 ;
        RECT 112.580 -2.825 112.880 4.105 ;
        RECT 113.890 -2.225 114.190 4.125 ;
        RECT 115.205 -2.195 115.500 4.630 ;
    END
  END s7
  PIN s7_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 122.070 4.180 122.450 4.560 ;
        RECT 118.995 3.685 121.620 4.095 ;
        RECT 121.180 1.245 124.255 1.520 ;
        RECT 121.195 -2.180 122.505 -1.860 ;
        RECT 119.005 -2.735 119.385 -2.355 ;
      LAYER Metal2 ;
        RECT 119.045 -2.825 119.345 4.115 ;
        RECT 121.255 -2.250 121.535 4.110 ;
        RECT 122.105 -2.250 122.405 4.570 ;
    END
  END s7_not
  PIN s1
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 114.990 122.735 115.370 123.115 ;
        RECT 112.315 122.310 114.055 122.600 ;
        RECT 113.670 117.715 124.075 118.050 ;
        RECT 113.640 116.395 115.420 116.685 ;
        RECT 112.370 115.780 112.750 116.160 ;
      LAYER Metal2 ;
        RECT 112.400 115.720 112.700 122.650 ;
        RECT 113.710 116.320 114.010 122.670 ;
        RECT 115.025 116.350 115.320 123.175 ;
    END
  END s1
  PIN s1_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 121.890 122.725 122.270 123.105 ;
        RECT 118.815 122.230 121.440 122.640 ;
        RECT 121.000 119.790 124.075 120.065 ;
        RECT 121.015 116.365 122.325 116.685 ;
        RECT 118.825 115.810 119.205 116.190 ;
      LAYER Metal2 ;
        RECT 118.865 115.720 119.165 122.660 ;
        RECT 121.075 116.295 121.355 122.655 ;
        RECT 121.925 116.295 122.225 123.115 ;
    END
  END s1_not
  PIN s6
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 115.170 23.855 115.550 24.235 ;
        RECT 112.495 23.430 114.235 23.720 ;
        RECT 113.850 18.835 124.255 19.170 ;
        RECT 113.820 17.515 115.600 17.805 ;
        RECT 112.550 16.900 112.930 17.280 ;
      LAYER Metal2 ;
        RECT 112.580 16.840 112.880 23.770 ;
        RECT 113.890 17.440 114.190 23.790 ;
        RECT 115.205 17.470 115.500 24.295 ;
    END
  END s6
  PIN s6_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 122.070 23.845 122.450 24.225 ;
        RECT 118.995 23.350 121.620 23.760 ;
        RECT 121.180 20.910 124.255 21.185 ;
        RECT 121.195 17.485 122.505 17.805 ;
        RECT 119.005 16.930 119.385 17.310 ;
      LAYER Metal2 ;
        RECT 119.045 16.840 119.345 23.780 ;
        RECT 121.255 17.415 121.535 23.775 ;
        RECT 122.105 17.415 122.405 24.235 ;
    END
  END s6_not
  PIN s0
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 115.190 142.460 115.570 142.840 ;
        RECT 112.515 142.035 114.255 142.325 ;
        RECT 113.870 137.440 124.275 137.775 ;
        RECT 113.840 136.120 115.620 136.410 ;
        RECT 112.570 135.505 112.950 135.885 ;
      LAYER Metal2 ;
        RECT 112.600 135.445 112.900 142.375 ;
        RECT 113.910 136.045 114.210 142.395 ;
        RECT 115.225 136.075 115.520 142.900 ;
    END
  END s0
  PIN s0_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 122.090 142.450 122.470 142.830 ;
        RECT 119.015 141.955 121.640 142.365 ;
        RECT 121.200 139.515 124.275 139.790 ;
        RECT 121.215 136.090 122.525 136.410 ;
        RECT 119.025 135.535 119.405 135.915 ;
      LAYER Metal2 ;
        RECT 119.065 135.445 119.365 142.385 ;
        RECT 121.275 136.020 121.555 142.380 ;
        RECT 122.125 136.020 122.425 142.840 ;
    END
  END s0_not
  PIN s5
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 115.170 43.825 115.550 44.205 ;
        RECT 112.495 43.400 114.235 43.690 ;
        RECT 113.850 38.805 124.255 39.140 ;
        RECT 113.820 37.485 115.600 37.775 ;
        RECT 112.550 36.870 112.930 37.250 ;
      LAYER Metal2 ;
        RECT 112.580 36.810 112.880 43.740 ;
        RECT 113.890 37.410 114.190 43.760 ;
        RECT 115.205 37.440 115.500 44.265 ;
    END
  END s5
  PIN s5_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 122.070 43.815 122.450 44.195 ;
        RECT 118.995 43.320 121.620 43.730 ;
        RECT 121.180 40.880 124.255 41.155 ;
        RECT 121.195 37.455 122.505 37.775 ;
        RECT 119.005 36.900 119.385 37.280 ;
      LAYER Metal2 ;
        RECT 119.045 36.810 119.345 43.750 ;
        RECT 121.255 37.385 121.535 43.745 ;
        RECT 122.105 37.385 122.405 44.205 ;
    END
  END s5_not
  PIN c15
    ANTENNADIFFAREA 2.734275 ;
    PORT
      LAYER Metal1 ;
        RECT 71.110 -173.655 71.490 -173.275 ;
        RECT 68.435 -174.080 70.175 -173.790 ;
        RECT 69.790 -178.675 80.195 -178.340 ;
        RECT 69.760 -179.995 71.540 -179.705 ;
        RECT 68.490 -180.610 68.870 -180.230 ;
      LAYER Metal2 ;
        RECT 68.520 -180.670 68.820 -173.740 ;
        RECT 69.830 -180.070 70.130 -173.720 ;
        RECT 71.145 -180.040 71.440 -173.215 ;
    END
  END c15
  PIN c15_not
    ANTENNADIFFAREA 2.560625 ;
    PORT
      LAYER Metal1 ;
        RECT 78.010 -173.665 78.390 -173.285 ;
        RECT 74.935 -174.175 77.635 -173.755 ;
        RECT 77.120 -176.600 80.195 -176.325 ;
        RECT 77.135 -180.025 78.445 -179.705 ;
        RECT 74.945 -180.580 75.325 -180.200 ;
      LAYER Metal2 ;
        RECT 74.985 -180.670 75.285 -173.730 ;
        RECT 77.195 -180.095 77.500 -173.735 ;
        RECT 78.045 -180.095 78.345 -173.275 ;
    END
  END c15_not
  PIN vdd
    ANTENNADIFFAREA 0.514800 ;
    PORT
      LAYER Nwell ;
        RECT 66.715 -176.525 82.175 -168.300 ;
      LAYER Metal1 ;
        RECT 66.715 -169.200 81.745 -168.300 ;
        RECT 80.995 -176.360 81.375 -169.200 ;
    END
  END vdd
  PIN vss
    ANTENNADIFFAREA 0.514800 ;
    PORT
      LAYER Pwell ;
        RECT 66.715 -184.225 82.175 -176.525 ;
      LAYER Metal1 ;
        RECT 66.715 -183.330 70.380 -183.320 ;
        RECT 80.995 -183.325 81.375 -177.495 ;
        RECT 80.625 -183.330 81.745 -183.325 ;
        RECT 66.715 -184.225 81.745 -183.330 ;
    END
  END vss
  PIN a15_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.405 -151.645 71.605 -151.265 ;
        RECT 70.405 -153.945 73.665 -153.565 ;
        RECT 71.070 -155.860 93.625 -155.520 ;
        RECT 94.735 -155.850 109.380 -155.550 ;
        RECT 70.385 -159.445 73.685 -159.065 ;
        RECT 97.760 -159.525 100.680 -159.225 ;
        RECT 104.225 -159.540 107.595 -159.240 ;
        RECT 70.385 -161.445 71.670 -161.065 ;
      LAYER Metal2 ;
        RECT 71.230 -162.175 71.545 -151.125 ;
        RECT 93.205 -155.930 93.625 -155.470 ;
        RECT 94.705 -155.935 95.125 -155.475 ;
        RECT 97.795 -159.575 98.095 -155.515 ;
        RECT 104.285 -159.590 104.565 -155.500 ;
        RECT 109.050 -155.980 109.355 -150.505 ;
      LAYER Metal3 ;
        RECT 109.005 -151.015 124.485 -150.560 ;
        RECT 93.175 -155.880 95.200 -155.495 ;
    END
  END a15_not_b
  PIN a15_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.930 -151.545 91.165 -151.165 ;
        RECT 87.905 -153.945 91.165 -153.565 ;
        RECT 95.335 -155.105 108.950 -154.805 ;
        RECT 96.530 -157.760 100.660 -157.460 ;
        RECT 103.035 -157.810 107.535 -157.500 ;
        RECT 89.790 -158.805 93.735 -158.470 ;
        RECT 87.885 -159.445 91.185 -159.065 ;
        RECT 89.700 -161.445 91.185 -161.065 ;
      LAYER Metal2 ;
        RECT 90.015 -161.690 90.330 -151.005 ;
        RECT 93.340 -158.820 93.720 -158.440 ;
        RECT 95.405 -158.845 95.715 -154.725 ;
        RECT 108.475 -155.150 108.770 -149.780 ;
      LAYER Metal3 ;
        RECT 108.475 -150.235 124.495 -149.825 ;
        RECT 93.340 -158.830 95.820 -158.430 ;
    END
  END a15_b
  PIN a14_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.405 -131.980 71.605 -131.600 ;
        RECT 70.405 -134.280 73.665 -133.900 ;
        RECT 71.070 -136.195 93.625 -135.855 ;
        RECT 94.735 -136.185 109.380 -135.885 ;
        RECT 70.385 -139.780 73.685 -139.400 ;
        RECT 97.760 -139.860 100.680 -139.560 ;
        RECT 104.225 -139.875 107.595 -139.575 ;
        RECT 70.385 -141.780 71.670 -141.400 ;
      LAYER Metal2 ;
        RECT 71.230 -142.510 71.545 -131.460 ;
        RECT 93.205 -136.265 93.625 -135.805 ;
        RECT 94.705 -136.270 95.125 -135.810 ;
        RECT 97.795 -139.910 98.095 -135.850 ;
        RECT 104.285 -139.925 104.565 -135.835 ;
        RECT 109.050 -136.315 109.355 -130.840 ;
      LAYER Metal3 ;
        RECT 109.005 -131.350 124.485 -130.895 ;
        RECT 93.175 -136.215 95.200 -135.830 ;
    END
  END a14_not_b
  PIN a14_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.930 -131.880 91.165 -131.500 ;
        RECT 87.905 -134.280 91.165 -133.900 ;
        RECT 95.335 -135.440 108.950 -135.140 ;
        RECT 96.530 -138.095 100.660 -137.795 ;
        RECT 103.035 -138.145 107.535 -137.835 ;
        RECT 89.790 -139.140 93.735 -138.805 ;
        RECT 87.885 -139.780 91.185 -139.400 ;
        RECT 89.700 -141.780 91.185 -141.400 ;
      LAYER Metal2 ;
        RECT 90.015 -142.025 90.330 -131.340 ;
        RECT 93.340 -139.155 93.720 -138.775 ;
        RECT 95.405 -139.180 95.715 -135.060 ;
        RECT 108.475 -135.485 108.770 -130.115 ;
      LAYER Metal3 ;
        RECT 108.475 -130.570 124.495 -130.160 ;
        RECT 93.340 -139.165 95.820 -138.765 ;
    END
  END a14_b
  PIN a13_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.405 -112.010 71.605 -111.630 ;
        RECT 70.405 -114.310 73.665 -113.930 ;
        RECT 71.070 -116.225 93.625 -115.885 ;
        RECT 94.735 -116.215 109.380 -115.915 ;
        RECT 70.385 -119.810 73.685 -119.430 ;
        RECT 97.760 -119.890 100.680 -119.590 ;
        RECT 104.225 -119.905 107.595 -119.605 ;
        RECT 70.385 -121.810 71.670 -121.430 ;
      LAYER Metal2 ;
        RECT 71.230 -122.540 71.545 -111.490 ;
        RECT 93.205 -116.295 93.625 -115.835 ;
        RECT 94.705 -116.300 95.125 -115.840 ;
        RECT 97.795 -119.940 98.095 -115.880 ;
        RECT 104.285 -119.955 104.565 -115.865 ;
        RECT 109.050 -116.345 109.355 -110.870 ;
      LAYER Metal3 ;
        RECT 109.005 -111.380 124.485 -110.925 ;
        RECT 93.175 -116.245 95.200 -115.860 ;
    END
  END a13_not_b
  PIN a13_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.930 -111.910 91.165 -111.530 ;
        RECT 87.905 -114.310 91.165 -113.930 ;
        RECT 95.335 -115.470 108.950 -115.170 ;
        RECT 96.530 -118.125 100.660 -117.825 ;
        RECT 103.035 -118.175 107.535 -117.865 ;
        RECT 89.790 -119.170 93.735 -118.835 ;
        RECT 87.885 -119.810 91.185 -119.430 ;
        RECT 89.700 -121.810 91.185 -121.430 ;
      LAYER Metal2 ;
        RECT 90.015 -122.055 90.330 -111.370 ;
        RECT 93.340 -119.185 93.720 -118.805 ;
        RECT 95.405 -119.210 95.715 -115.090 ;
        RECT 108.475 -115.515 108.770 -110.145 ;
      LAYER Metal3 ;
        RECT 108.475 -110.600 124.495 -110.190 ;
        RECT 93.340 -119.195 95.820 -118.795 ;
    END
  END a13_b
  PIN a12_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.300 -92.295 71.500 -91.915 ;
        RECT 70.300 -94.595 73.560 -94.215 ;
        RECT 70.965 -96.510 93.520 -96.170 ;
        RECT 94.630 -96.500 109.275 -96.200 ;
        RECT 70.280 -100.095 73.580 -99.715 ;
        RECT 97.655 -100.175 100.575 -99.875 ;
        RECT 104.120 -100.190 107.490 -99.890 ;
        RECT 70.280 -102.095 71.565 -101.715 ;
      LAYER Metal2 ;
        RECT 71.125 -102.825 71.440 -91.775 ;
        RECT 93.100 -96.580 93.520 -96.120 ;
        RECT 94.600 -96.585 95.020 -96.125 ;
        RECT 97.690 -100.225 97.990 -96.165 ;
        RECT 104.180 -100.240 104.460 -96.150 ;
        RECT 108.945 -96.630 109.250 -91.155 ;
      LAYER Metal3 ;
        RECT 108.900 -91.665 124.380 -91.210 ;
        RECT 93.070 -96.530 95.095 -96.145 ;
    END
  END a12_not_b
  PIN a12_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.825 -92.195 91.060 -91.815 ;
        RECT 87.800 -94.595 91.060 -94.215 ;
        RECT 95.230 -95.755 108.845 -95.455 ;
        RECT 96.425 -98.410 100.555 -98.110 ;
        RECT 102.930 -98.460 107.430 -98.150 ;
        RECT 89.685 -99.455 93.630 -99.120 ;
        RECT 87.780 -100.095 91.080 -99.715 ;
        RECT 89.595 -102.095 91.080 -101.715 ;
      LAYER Metal2 ;
        RECT 89.910 -102.340 90.225 -91.655 ;
        RECT 93.235 -99.470 93.615 -99.090 ;
        RECT 95.300 -99.495 95.610 -95.375 ;
        RECT 108.370 -95.800 108.665 -90.430 ;
      LAYER Metal3 ;
        RECT 108.370 -90.885 124.390 -90.475 ;
        RECT 93.235 -99.480 95.715 -99.080 ;
    END
  END a12_b
  PIN a11_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.380 -72.540 71.580 -72.160 ;
        RECT 70.380 -74.840 73.640 -74.460 ;
        RECT 71.045 -76.755 93.600 -76.415 ;
        RECT 94.710 -76.745 109.355 -76.445 ;
        RECT 70.360 -80.340 73.660 -79.960 ;
        RECT 97.735 -80.420 100.655 -80.120 ;
        RECT 104.200 -80.435 107.570 -80.135 ;
        RECT 70.360 -82.340 71.645 -81.960 ;
      LAYER Metal2 ;
        RECT 71.205 -83.070 71.520 -72.020 ;
        RECT 93.180 -76.825 93.600 -76.365 ;
        RECT 94.680 -76.830 95.100 -76.370 ;
        RECT 97.770 -80.470 98.070 -76.410 ;
        RECT 104.260 -80.485 104.540 -76.395 ;
        RECT 109.025 -76.875 109.330 -71.400 ;
      LAYER Metal3 ;
        RECT 108.980 -71.910 124.460 -71.455 ;
        RECT 93.150 -76.775 95.175 -76.390 ;
    END
  END a11_not_b
  PIN a11_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.905 -72.440 91.140 -72.060 ;
        RECT 87.880 -74.840 91.140 -74.460 ;
        RECT 95.310 -76.000 108.925 -75.700 ;
        RECT 96.505 -78.655 100.635 -78.355 ;
        RECT 103.010 -78.705 107.510 -78.395 ;
        RECT 89.765 -79.700 93.710 -79.365 ;
        RECT 87.860 -80.340 91.160 -79.960 ;
        RECT 89.675 -82.340 91.160 -81.960 ;
      LAYER Metal2 ;
        RECT 89.990 -82.585 90.305 -71.900 ;
        RECT 93.315 -79.715 93.695 -79.335 ;
        RECT 95.380 -79.740 95.690 -75.620 ;
        RECT 108.450 -76.045 108.745 -70.675 ;
      LAYER Metal3 ;
        RECT 108.450 -71.130 124.470 -70.720 ;
        RECT 93.315 -79.725 95.795 -79.325 ;
    END
  END a11_b
  PIN a10_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.380 -52.745 71.580 -52.365 ;
        RECT 70.380 -55.045 73.640 -54.665 ;
        RECT 71.045 -56.960 93.600 -56.620 ;
        RECT 94.710 -56.950 109.355 -56.650 ;
        RECT 70.360 -60.545 73.660 -60.165 ;
        RECT 97.735 -60.625 100.655 -60.325 ;
        RECT 104.200 -60.640 107.570 -60.340 ;
        RECT 70.360 -62.545 71.645 -62.165 ;
      LAYER Metal2 ;
        RECT 71.205 -63.275 71.520 -52.225 ;
        RECT 93.180 -57.030 93.600 -56.570 ;
        RECT 94.680 -57.035 95.100 -56.575 ;
        RECT 97.770 -60.675 98.070 -56.615 ;
        RECT 104.260 -60.690 104.540 -56.600 ;
        RECT 109.025 -57.080 109.330 -51.605 ;
      LAYER Metal3 ;
        RECT 108.980 -52.115 124.460 -51.660 ;
        RECT 93.150 -56.980 95.175 -56.595 ;
    END
  END a10_not_b
  PIN a10_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.905 -52.645 91.140 -52.265 ;
        RECT 87.880 -55.045 91.140 -54.665 ;
        RECT 95.310 -56.205 108.925 -55.905 ;
        RECT 96.505 -58.860 100.635 -58.560 ;
        RECT 103.010 -58.910 107.510 -58.600 ;
        RECT 89.765 -59.905 93.710 -59.570 ;
        RECT 87.860 -60.545 91.160 -60.165 ;
        RECT 89.675 -62.545 91.160 -62.165 ;
      LAYER Metal2 ;
        RECT 89.990 -62.790 90.305 -52.105 ;
        RECT 93.315 -59.920 93.695 -59.540 ;
        RECT 95.380 -59.945 95.690 -55.825 ;
        RECT 108.450 -56.250 108.745 -50.880 ;
      LAYER Metal3 ;
        RECT 108.450 -51.335 124.470 -50.925 ;
        RECT 93.315 -59.930 95.795 -59.530 ;
    END
  END a10_b
  PIN a9_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.225 -33.100 71.425 -32.720 ;
        RECT 70.225 -35.400 73.485 -35.020 ;
        RECT 70.890 -37.315 93.445 -36.975 ;
        RECT 94.555 -37.305 109.200 -37.005 ;
        RECT 70.205 -40.900 73.505 -40.520 ;
        RECT 97.580 -40.980 100.500 -40.680 ;
        RECT 104.045 -40.995 107.415 -40.695 ;
        RECT 70.205 -42.900 71.490 -42.520 ;
      LAYER Metal2 ;
        RECT 71.050 -43.630 71.365 -32.580 ;
        RECT 93.025 -37.385 93.445 -36.925 ;
        RECT 94.525 -37.390 94.945 -36.930 ;
        RECT 97.615 -41.030 97.915 -36.970 ;
        RECT 104.105 -41.045 104.385 -36.955 ;
        RECT 108.870 -37.435 109.175 -31.960 ;
      LAYER Metal3 ;
        RECT 108.825 -32.470 124.305 -32.015 ;
        RECT 92.995 -37.335 95.020 -36.950 ;
    END
  END a9_not_b
  PIN a9_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.750 -33.000 90.985 -32.620 ;
        RECT 87.725 -35.400 90.985 -35.020 ;
        RECT 95.155 -36.560 108.770 -36.260 ;
        RECT 96.350 -39.215 100.480 -38.915 ;
        RECT 102.855 -39.265 107.355 -38.955 ;
        RECT 89.610 -40.260 93.555 -39.925 ;
        RECT 87.705 -40.900 91.005 -40.520 ;
        RECT 89.520 -42.900 91.005 -42.520 ;
      LAYER Metal2 ;
        RECT 89.835 -43.145 90.150 -32.460 ;
        RECT 93.160 -40.275 93.540 -39.895 ;
        RECT 95.225 -40.300 95.535 -36.180 ;
        RECT 108.295 -36.605 108.590 -31.235 ;
      LAYER Metal3 ;
        RECT 108.295 -31.690 124.315 -31.280 ;
        RECT 93.160 -40.285 95.640 -39.885 ;
    END
  END a9_b
  PIN a8_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.425 -13.375 71.625 -12.995 ;
        RECT 70.425 -15.675 73.685 -15.295 ;
        RECT 71.090 -17.590 93.645 -17.250 ;
        RECT 94.755 -17.580 109.400 -17.280 ;
        RECT 70.405 -21.175 73.705 -20.795 ;
        RECT 97.780 -21.255 100.700 -20.955 ;
        RECT 104.245 -21.270 107.615 -20.970 ;
        RECT 70.405 -23.175 71.690 -22.795 ;
      LAYER Metal2 ;
        RECT 71.250 -23.905 71.565 -12.855 ;
        RECT 93.225 -17.660 93.645 -17.200 ;
        RECT 94.725 -17.665 95.145 -17.205 ;
        RECT 97.815 -21.305 98.115 -17.245 ;
        RECT 104.305 -21.320 104.585 -17.230 ;
        RECT 109.070 -17.710 109.375 -12.235 ;
      LAYER Metal3 ;
        RECT 109.025 -12.745 124.505 -12.290 ;
        RECT 93.195 -17.610 95.220 -17.225 ;
    END
  END a8_not_b
  PIN a8_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.950 -13.275 91.185 -12.895 ;
        RECT 87.925 -15.675 91.185 -15.295 ;
        RECT 95.355 -16.835 108.970 -16.535 ;
        RECT 96.550 -19.490 100.680 -19.190 ;
        RECT 103.055 -19.540 107.555 -19.230 ;
        RECT 89.810 -20.535 93.755 -20.200 ;
        RECT 87.905 -21.175 91.205 -20.795 ;
        RECT 89.720 -23.175 91.205 -22.795 ;
      LAYER Metal2 ;
        RECT 90.035 -23.420 90.350 -12.735 ;
        RECT 93.360 -20.550 93.740 -20.170 ;
        RECT 95.425 -20.575 95.735 -16.455 ;
        RECT 108.495 -16.880 108.790 -11.510 ;
      LAYER Metal3 ;
        RECT 108.495 -11.965 124.515 -11.555 ;
        RECT 93.360 -20.560 95.840 -20.160 ;
    END
  END a8_b
  PIN a7_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.385 6.465 71.585 6.845 ;
        RECT 70.385 4.165 73.645 4.545 ;
        RECT 71.050 2.250 93.605 2.590 ;
        RECT 94.715 2.260 109.360 2.560 ;
        RECT 70.365 -1.335 73.665 -0.955 ;
        RECT 97.740 -1.415 100.660 -1.115 ;
        RECT 104.205 -1.430 107.575 -1.130 ;
        RECT 70.365 -3.335 71.650 -2.955 ;
      LAYER Metal2 ;
        RECT 71.210 -4.065 71.525 6.985 ;
        RECT 93.185 2.180 93.605 2.640 ;
        RECT 94.685 2.175 95.105 2.635 ;
        RECT 97.775 -1.465 98.075 2.595 ;
        RECT 104.265 -1.480 104.545 2.610 ;
        RECT 109.030 2.130 109.335 7.605 ;
      LAYER Metal3 ;
        RECT 108.985 7.095 124.465 7.550 ;
        RECT 93.155 2.230 95.180 2.615 ;
    END
  END a7_not_b
  PIN a7_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.910 6.565 91.145 6.945 ;
        RECT 87.885 4.165 91.145 4.545 ;
        RECT 95.315 3.005 108.930 3.305 ;
        RECT 96.510 0.350 100.640 0.650 ;
        RECT 103.015 0.300 107.515 0.610 ;
        RECT 89.770 -0.695 93.715 -0.360 ;
        RECT 87.865 -1.335 91.165 -0.955 ;
        RECT 89.680 -3.335 91.165 -2.955 ;
      LAYER Metal2 ;
        RECT 89.995 -3.580 90.310 7.105 ;
        RECT 93.320 -0.710 93.700 -0.330 ;
        RECT 95.385 -0.735 95.695 3.385 ;
        RECT 108.455 2.960 108.750 8.330 ;
      LAYER Metal3 ;
        RECT 108.455 7.875 124.475 8.285 ;
        RECT 93.320 -0.720 95.800 -0.320 ;
    END
  END a7_b
  PIN a6_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.385 26.130 71.585 26.510 ;
        RECT 70.385 23.830 73.645 24.210 ;
        RECT 71.050 21.915 93.605 22.255 ;
        RECT 94.715 21.925 109.360 22.225 ;
        RECT 70.365 18.330 73.665 18.710 ;
        RECT 97.740 18.250 100.660 18.550 ;
        RECT 104.205 18.235 107.575 18.535 ;
        RECT 70.365 16.330 71.650 16.710 ;
      LAYER Metal2 ;
        RECT 71.210 15.600 71.525 26.650 ;
        RECT 93.185 21.845 93.605 22.305 ;
        RECT 94.685 21.840 95.105 22.300 ;
        RECT 97.775 18.200 98.075 22.260 ;
        RECT 104.265 18.185 104.545 22.275 ;
        RECT 109.030 21.795 109.335 27.270 ;
      LAYER Metal3 ;
        RECT 108.985 26.760 124.465 27.215 ;
        RECT 93.155 21.895 95.180 22.280 ;
    END
  END a6_not_b
  PIN a6_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.910 26.230 91.145 26.610 ;
        RECT 87.885 23.830 91.145 24.210 ;
        RECT 95.315 22.670 108.930 22.970 ;
        RECT 96.510 20.015 100.640 20.315 ;
        RECT 103.015 19.965 107.515 20.275 ;
        RECT 89.770 18.970 93.715 19.305 ;
        RECT 87.865 18.330 91.165 18.710 ;
        RECT 89.680 16.330 91.165 16.710 ;
      LAYER Metal2 ;
        RECT 89.995 16.085 90.310 26.770 ;
        RECT 93.320 18.955 93.700 19.335 ;
        RECT 95.385 18.930 95.695 23.050 ;
        RECT 108.455 22.625 108.750 27.995 ;
      LAYER Metal3 ;
        RECT 108.455 27.540 124.475 27.950 ;
        RECT 93.320 18.945 95.800 19.345 ;
    END
  END a6_b
  PIN a5_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.385 46.100 71.585 46.480 ;
        RECT 70.385 43.800 73.645 44.180 ;
        RECT 71.050 41.885 93.605 42.225 ;
        RECT 94.715 41.895 109.360 42.195 ;
        RECT 70.365 38.300 73.665 38.680 ;
        RECT 97.740 38.220 100.660 38.520 ;
        RECT 104.205 38.205 107.575 38.505 ;
        RECT 70.365 36.300 71.650 36.680 ;
      LAYER Metal2 ;
        RECT 71.210 35.570 71.525 46.620 ;
        RECT 93.185 41.815 93.605 42.275 ;
        RECT 94.685 41.810 95.105 42.270 ;
        RECT 97.775 38.170 98.075 42.230 ;
        RECT 104.265 38.155 104.545 42.245 ;
        RECT 109.030 41.765 109.335 47.240 ;
      LAYER Metal3 ;
        RECT 108.985 46.730 124.465 47.185 ;
        RECT 93.155 41.865 95.180 42.250 ;
    END
  END a5_not_b
  PIN a5_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.910 46.200 91.145 46.580 ;
        RECT 87.885 43.800 91.145 44.180 ;
        RECT 95.315 42.640 108.930 42.940 ;
        RECT 96.510 39.985 100.640 40.285 ;
        RECT 103.015 39.935 107.515 40.245 ;
        RECT 89.770 38.940 93.715 39.275 ;
        RECT 87.865 38.300 91.165 38.680 ;
        RECT 89.680 36.300 91.165 36.680 ;
      LAYER Metal2 ;
        RECT 89.995 36.055 90.310 46.740 ;
        RECT 93.320 38.925 93.700 39.305 ;
        RECT 95.385 38.900 95.695 43.020 ;
        RECT 108.455 42.595 108.750 47.965 ;
      LAYER Metal3 ;
        RECT 108.455 47.510 124.475 47.920 ;
        RECT 93.320 38.915 95.800 39.315 ;
    END
  END a5_b
  PIN a4_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.280 65.815 71.480 66.195 ;
        RECT 70.280 63.515 73.540 63.895 ;
        RECT 70.945 61.600 93.500 61.940 ;
        RECT 94.610 61.610 109.255 61.910 ;
        RECT 70.260 58.015 73.560 58.395 ;
        RECT 97.635 57.935 100.555 58.235 ;
        RECT 104.100 57.920 107.470 58.220 ;
        RECT 70.260 56.015 71.545 56.395 ;
      LAYER Metal2 ;
        RECT 71.105 55.285 71.420 66.335 ;
        RECT 93.080 61.530 93.500 61.990 ;
        RECT 94.580 61.525 95.000 61.985 ;
        RECT 97.670 57.885 97.970 61.945 ;
        RECT 104.160 57.870 104.440 61.960 ;
        RECT 108.925 61.480 109.230 66.955 ;
      LAYER Metal3 ;
        RECT 108.880 66.445 124.360 66.900 ;
        RECT 93.050 61.580 95.075 61.965 ;
    END
  END a4_not_b
  PIN a4_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.805 65.915 91.040 66.295 ;
        RECT 87.780 63.515 91.040 63.895 ;
        RECT 95.210 62.355 108.825 62.655 ;
        RECT 96.405 59.700 100.535 60.000 ;
        RECT 102.910 59.650 107.410 59.960 ;
        RECT 89.665 58.655 93.610 58.990 ;
        RECT 87.760 58.015 91.060 58.395 ;
        RECT 89.575 56.015 91.060 56.395 ;
      LAYER Metal2 ;
        RECT 89.890 55.770 90.205 66.455 ;
        RECT 93.215 58.640 93.595 59.020 ;
        RECT 95.280 58.615 95.590 62.735 ;
        RECT 108.350 62.310 108.645 67.680 ;
      LAYER Metal3 ;
        RECT 108.350 67.225 124.370 67.635 ;
        RECT 93.215 58.630 95.695 59.030 ;
    END
  END a4_b
  PIN a3_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.360 85.570 71.560 85.950 ;
        RECT 70.360 83.270 73.620 83.650 ;
        RECT 71.025 81.355 93.580 81.695 ;
        RECT 94.690 81.365 109.335 81.665 ;
        RECT 70.340 77.770 73.640 78.150 ;
        RECT 97.715 77.690 100.635 77.990 ;
        RECT 104.180 77.675 107.550 77.975 ;
        RECT 70.340 75.770 71.625 76.150 ;
      LAYER Metal2 ;
        RECT 71.185 75.040 71.500 86.090 ;
        RECT 93.160 81.285 93.580 81.745 ;
        RECT 94.660 81.280 95.080 81.740 ;
        RECT 97.750 77.640 98.050 81.700 ;
        RECT 104.240 77.625 104.520 81.715 ;
        RECT 109.005 81.235 109.310 86.710 ;
      LAYER Metal3 ;
        RECT 108.960 86.200 124.440 86.655 ;
        RECT 93.130 81.335 95.155 81.720 ;
    END
  END a3_not_b
  PIN a3_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.885 85.670 91.120 86.050 ;
        RECT 87.860 83.270 91.120 83.650 ;
        RECT 95.290 82.110 108.905 82.410 ;
        RECT 96.485 79.455 100.615 79.755 ;
        RECT 102.990 79.405 107.490 79.715 ;
        RECT 89.745 78.410 93.690 78.745 ;
        RECT 87.840 77.770 91.140 78.150 ;
        RECT 89.655 75.770 91.140 76.150 ;
      LAYER Metal2 ;
        RECT 89.970 75.525 90.285 86.210 ;
        RECT 93.295 78.395 93.675 78.775 ;
        RECT 95.360 78.370 95.670 82.490 ;
        RECT 108.430 82.065 108.725 87.435 ;
      LAYER Metal3 ;
        RECT 108.430 86.980 124.450 87.390 ;
        RECT 93.295 78.385 95.775 78.785 ;
    END
  END a3_b
  PIN a2_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.360 105.365 71.560 105.745 ;
        RECT 70.360 103.065 73.620 103.445 ;
        RECT 71.025 101.150 93.580 101.490 ;
        RECT 94.690 101.160 109.335 101.460 ;
        RECT 70.340 97.565 73.640 97.945 ;
        RECT 97.715 97.485 100.635 97.785 ;
        RECT 104.180 97.470 107.550 97.770 ;
        RECT 70.340 95.565 71.625 95.945 ;
      LAYER Metal2 ;
        RECT 71.185 94.835 71.500 105.885 ;
        RECT 93.160 101.080 93.580 101.540 ;
        RECT 94.660 101.075 95.080 101.535 ;
        RECT 97.750 97.435 98.050 101.495 ;
        RECT 104.240 97.420 104.520 101.510 ;
        RECT 109.005 101.030 109.310 106.505 ;
      LAYER Metal3 ;
        RECT 108.960 105.995 124.440 106.450 ;
        RECT 93.130 101.130 95.155 101.515 ;
    END
  END a2_not_b
  PIN a2_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.885 105.465 91.120 105.845 ;
        RECT 87.860 103.065 91.120 103.445 ;
        RECT 95.290 101.905 108.905 102.205 ;
        RECT 96.485 99.250 100.615 99.550 ;
        RECT 102.990 99.200 107.490 99.510 ;
        RECT 89.745 98.205 93.690 98.540 ;
        RECT 87.840 97.565 91.140 97.945 ;
        RECT 89.655 95.565 91.140 95.945 ;
      LAYER Metal2 ;
        RECT 89.970 95.320 90.285 106.005 ;
        RECT 93.295 98.190 93.675 98.570 ;
        RECT 95.360 98.165 95.670 102.285 ;
        RECT 108.430 101.860 108.725 107.230 ;
      LAYER Metal3 ;
        RECT 108.430 106.775 124.450 107.185 ;
        RECT 93.295 98.180 95.775 98.580 ;
    END
  END a2_b
  PIN a1_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.205 125.010 71.405 125.390 ;
        RECT 70.205 122.710 73.465 123.090 ;
        RECT 70.870 120.795 93.425 121.135 ;
        RECT 94.535 120.805 109.180 121.105 ;
        RECT 70.185 117.210 73.485 117.590 ;
        RECT 97.560 117.130 100.480 117.430 ;
        RECT 104.025 117.115 107.395 117.415 ;
        RECT 70.185 115.210 71.470 115.590 ;
      LAYER Metal2 ;
        RECT 71.030 114.480 71.345 125.530 ;
        RECT 93.005 120.725 93.425 121.185 ;
        RECT 94.505 120.720 94.925 121.180 ;
        RECT 97.595 117.080 97.895 121.140 ;
        RECT 104.085 117.065 104.365 121.155 ;
        RECT 108.850 120.675 109.155 126.150 ;
      LAYER Metal3 ;
        RECT 108.805 125.640 124.285 126.095 ;
        RECT 92.975 120.775 95.000 121.160 ;
    END
  END a1_not_b
  PIN a1_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.730 125.110 90.965 125.490 ;
        RECT 87.705 122.710 90.965 123.090 ;
        RECT 95.135 121.550 108.750 121.850 ;
        RECT 96.330 118.895 100.460 119.195 ;
        RECT 102.835 118.845 107.335 119.155 ;
        RECT 89.590 117.850 93.535 118.185 ;
        RECT 87.685 117.210 90.985 117.590 ;
        RECT 89.500 115.210 90.985 115.590 ;
      LAYER Metal2 ;
        RECT 89.815 114.965 90.130 125.650 ;
        RECT 93.140 117.835 93.520 118.215 ;
        RECT 95.205 117.810 95.515 121.930 ;
        RECT 108.275 121.505 108.570 126.875 ;
      LAYER Metal3 ;
        RECT 108.275 126.420 124.295 126.830 ;
        RECT 93.140 117.825 95.620 118.225 ;
    END
  END a1_b
  PIN a0_not_b
    ANTENNAGATEAREA 2.775000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 70.405 144.735 71.605 145.115 ;
        RECT 70.405 142.435 73.665 142.815 ;
        RECT 71.070 140.520 93.625 140.860 ;
        RECT 94.735 140.530 109.380 140.830 ;
        RECT 70.385 136.935 73.685 137.315 ;
        RECT 97.760 136.855 100.680 137.155 ;
        RECT 104.225 136.840 107.595 137.140 ;
        RECT 70.385 134.935 71.670 135.315 ;
      LAYER Metal2 ;
        RECT 71.230 134.205 71.545 145.255 ;
        RECT 93.205 140.450 93.625 140.910 ;
        RECT 94.705 140.445 95.125 140.905 ;
        RECT 97.795 136.805 98.095 140.865 ;
        RECT 104.285 136.790 104.565 140.880 ;
        RECT 109.050 140.400 109.355 145.875 ;
      LAYER Metal3 ;
        RECT 109.005 145.365 124.485 145.820 ;
        RECT 93.175 140.500 95.200 140.885 ;
    END
  END a0_not_b
  PIN a0_b
    ANTENNAGATEAREA 2.739250 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 89.930 144.835 91.165 145.215 ;
        RECT 87.905 142.435 91.165 142.815 ;
        RECT 95.335 141.275 108.950 141.575 ;
        RECT 96.530 138.620 100.660 138.920 ;
        RECT 103.035 138.570 107.535 138.880 ;
        RECT 89.790 137.575 93.735 137.910 ;
        RECT 87.885 136.935 91.185 137.315 ;
        RECT 89.700 134.935 91.185 135.315 ;
      LAYER Metal2 ;
        RECT 90.015 134.690 90.330 145.375 ;
        RECT 93.340 137.560 93.720 137.940 ;
        RECT 95.405 137.535 95.715 141.655 ;
        RECT 108.475 141.230 108.770 146.600 ;
      LAYER Metal3 ;
        RECT 108.475 146.145 124.495 146.555 ;
        RECT 93.340 137.550 95.820 137.950 ;
    END
  END a0_b
  PIN b15_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -2.270 -153.670 1.105 -153.270 ;
        RECT 9.510 -154.320 9.890 -153.940 ;
        RECT -2.960 -157.175 1.165 -156.905 ;
        RECT 0.740 -158.350 7.130 -158.060 ;
        RECT -2.280 -160.265 -1.900 -159.885 ;
        RECT 6.720 -160.990 9.900 -160.670 ;
      LAYER Metal2 ;
        RECT -2.950 -157.245 -2.570 -156.865 ;
        RECT -2.235 -160.320 -1.935 -153.280 ;
        RECT 0.790 -158.450 1.110 -153.290 ;
        RECT 6.800 -161.050 7.080 -158.015 ;
        RECT 9.550 -161.095 9.850 -153.940 ;
      LAYER Metal3 ;
        RECT -5.360 -157.180 -2.565 -156.885 ;
    END
  END b15_not
  PIN b15
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.190 -153.870 4.570 -153.490 ;
        RECT 2.590 -154.385 3.790 -154.095 ;
        RECT -2.940 -156.555 3.785 -156.255 ;
        RECT 3.380 -160.160 4.570 -159.875 ;
        RECT 2.600 -160.825 2.980 -160.445 ;
      LAYER Metal2 ;
        RECT -2.915 -156.575 -2.535 -156.195 ;
        RECT 2.640 -160.835 2.940 -154.025 ;
        RECT 3.430 -160.240 3.740 -154.050 ;
        RECT 4.225 -160.310 4.525 -153.480 ;
      LAYER Metal3 ;
        RECT -5.395 -156.550 -2.520 -156.255 ;
    END
  END b15
  PIN a15_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.510 -151.635 30.965 -151.255 ;
        RECT 29.670 -153.935 30.965 -153.555 ;
        RECT 43.155 -153.935 44.465 -153.555 ;
        RECT 28.000 -155.260 44.010 -154.885 ;
        RECT -2.960 -155.840 10.600 -155.540 ;
        RECT 12.505 -155.840 30.925 -155.540 ;
        RECT -0.495 -159.515 2.425 -159.215 ;
        RECT 5.970 -159.530 9.340 -159.230 ;
        RECT 14.965 -159.515 17.885 -159.215 ;
        RECT 21.430 -159.530 24.800 -159.230 ;
        RECT 29.680 -159.435 30.985 -159.055 ;
        RECT 43.020 -159.435 44.485 -159.055 ;
        RECT 29.495 -161.435 30.985 -161.055 ;
      LAYER Metal2 ;
        RECT -2.960 -155.890 -2.580 -155.510 ;
        RECT -0.460 -159.565 -0.160 -155.505 ;
        RECT 6.030 -159.580 6.310 -155.490 ;
        RECT 10.220 -155.890 10.600 -155.510 ;
        RECT 12.490 -155.890 12.870 -155.485 ;
        RECT 15.000 -159.565 15.300 -155.505 ;
        RECT 21.490 -159.580 21.770 -155.490 ;
        RECT 29.800 -161.490 30.155 -151.185 ;
        RECT 30.465 -155.885 30.810 -154.830 ;
        RECT 43.310 -159.715 43.640 -153.520 ;
      LAYER Metal3 ;
        RECT -5.400 -155.835 -2.555 -155.540 ;
        RECT 10.165 -155.860 12.905 -155.530 ;
    END
  END a15_not_f
  PIN a15_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.205 -151.535 54.485 -151.155 ;
        RECT 39.705 -153.935 40.890 -153.555 ;
        RECT 53.205 -153.935 54.220 -153.555 ;
        RECT -2.955 -155.095 10.610 -154.780 ;
        RECT 12.500 -155.095 26.325 -154.795 ;
        RECT 28.000 -156.615 54.230 -156.225 ;
        RECT -1.725 -157.750 2.405 -157.450 ;
        RECT 4.780 -157.800 9.280 -157.490 ;
        RECT 13.735 -157.750 17.865 -157.450 ;
        RECT 20.240 -157.800 24.740 -157.490 ;
        RECT 39.685 -159.435 41.045 -159.055 ;
        RECT 53.185 -159.435 54.365 -159.055 ;
        RECT 53.185 -161.435 54.260 -161.055 ;
      LAYER Metal2 ;
        RECT -2.950 -155.140 -2.570 -154.760 ;
        RECT 10.215 -155.140 10.595 -154.760 ;
        RECT 12.485 -155.140 12.865 -154.735 ;
        RECT 25.950 -155.140 26.310 -153.310 ;
        RECT 28.130 -156.660 28.545 -153.310 ;
        RECT 40.325 -153.570 40.635 -153.540 ;
        RECT 40.325 -159.670 40.640 -153.570 ;
        RECT 53.825 -161.665 54.155 -150.970 ;
      LAYER Metal3 ;
        RECT 25.895 -153.695 28.600 -153.355 ;
        RECT -5.360 -155.100 -2.535 -154.795 ;
        RECT 10.160 -155.110 12.905 -154.780 ;
    END
  END a15_f
  PIN b14_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -2.240 -133.875 1.135 -133.475 ;
        RECT 9.540 -134.525 9.920 -134.145 ;
        RECT -2.930 -137.380 1.195 -137.110 ;
        RECT 0.770 -138.555 7.160 -138.265 ;
        RECT -2.250 -140.470 -1.870 -140.090 ;
        RECT 6.750 -141.195 9.930 -140.875 ;
      LAYER Metal2 ;
        RECT -2.920 -137.450 -2.540 -137.070 ;
        RECT -2.205 -140.525 -1.905 -133.485 ;
        RECT 0.820 -138.655 1.140 -133.495 ;
        RECT 6.830 -141.255 7.110 -138.220 ;
        RECT 9.580 -141.300 9.880 -134.145 ;
      LAYER Metal3 ;
        RECT -5.330 -137.385 -2.535 -137.090 ;
    END
  END b14_not
  PIN b14
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.220 -134.075 4.600 -133.695 ;
        RECT 2.620 -134.590 3.820 -134.300 ;
        RECT -2.910 -136.760 3.815 -136.460 ;
        RECT 3.410 -140.365 4.600 -140.080 ;
        RECT 2.630 -141.030 3.010 -140.650 ;
      LAYER Metal2 ;
        RECT -2.885 -136.780 -2.505 -136.400 ;
        RECT 2.670 -141.040 2.970 -134.230 ;
        RECT 3.460 -140.445 3.770 -134.255 ;
        RECT 4.255 -140.515 4.555 -133.685 ;
      LAYER Metal3 ;
        RECT -5.365 -136.755 -2.490 -136.460 ;
    END
  END b14
  PIN a14_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.540 -131.840 30.995 -131.460 ;
        RECT 29.700 -134.140 30.995 -133.760 ;
        RECT 43.185 -134.140 44.495 -133.760 ;
        RECT 28.030 -135.465 44.040 -135.090 ;
        RECT -2.930 -136.045 10.630 -135.745 ;
        RECT 12.535 -136.045 30.955 -135.745 ;
        RECT -0.465 -139.720 2.455 -139.420 ;
        RECT 6.000 -139.735 9.370 -139.435 ;
        RECT 14.995 -139.720 17.915 -139.420 ;
        RECT 21.460 -139.735 24.830 -139.435 ;
        RECT 29.710 -139.640 31.015 -139.260 ;
        RECT 43.050 -139.640 44.515 -139.260 ;
        RECT 29.525 -141.640 31.015 -141.260 ;
      LAYER Metal2 ;
        RECT -2.930 -136.095 -2.550 -135.715 ;
        RECT -0.430 -139.770 -0.130 -135.710 ;
        RECT 6.060 -139.785 6.340 -135.695 ;
        RECT 10.250 -136.095 10.630 -135.715 ;
        RECT 12.520 -136.095 12.900 -135.690 ;
        RECT 15.030 -139.770 15.330 -135.710 ;
        RECT 21.520 -139.785 21.800 -135.695 ;
        RECT 29.830 -141.695 30.185 -131.390 ;
        RECT 30.495 -136.090 30.840 -135.035 ;
        RECT 43.340 -139.920 43.670 -133.725 ;
      LAYER Metal3 ;
        RECT -5.370 -136.040 -2.525 -135.745 ;
        RECT 10.195 -136.065 12.935 -135.735 ;
    END
  END a14_not_f
  PIN a14_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.235 -131.740 54.515 -131.360 ;
        RECT 39.735 -134.140 40.920 -133.760 ;
        RECT 53.235 -134.140 54.250 -133.760 ;
        RECT -2.925 -135.300 10.640 -134.985 ;
        RECT 12.530 -135.300 26.355 -135.000 ;
        RECT 28.030 -136.820 54.260 -136.430 ;
        RECT -1.695 -137.955 2.435 -137.655 ;
        RECT 4.810 -138.005 9.310 -137.695 ;
        RECT 13.765 -137.955 17.895 -137.655 ;
        RECT 20.270 -138.005 24.770 -137.695 ;
        RECT 39.715 -139.640 41.075 -139.260 ;
        RECT 53.215 -139.640 54.395 -139.260 ;
        RECT 53.215 -141.640 54.290 -141.260 ;
      LAYER Metal2 ;
        RECT -2.920 -135.345 -2.540 -134.965 ;
        RECT 10.245 -135.345 10.625 -134.965 ;
        RECT 12.515 -135.345 12.895 -134.940 ;
        RECT 25.980 -135.345 26.340 -133.515 ;
        RECT 28.160 -136.865 28.575 -133.515 ;
        RECT 40.355 -133.775 40.665 -133.745 ;
        RECT 40.355 -139.875 40.670 -133.775 ;
        RECT 53.855 -141.870 54.185 -131.175 ;
      LAYER Metal3 ;
        RECT 25.925 -133.900 28.630 -133.560 ;
        RECT -5.330 -135.305 -2.505 -135.000 ;
        RECT 10.190 -135.315 12.935 -134.985 ;
    END
  END a14_f
  PIN b13_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -2.190 -114.065 1.185 -113.665 ;
        RECT 9.590 -114.715 9.970 -114.335 ;
        RECT -2.880 -117.570 1.245 -117.300 ;
        RECT 0.820 -118.745 7.210 -118.455 ;
        RECT -2.200 -120.660 -1.820 -120.280 ;
        RECT 6.800 -121.385 9.980 -121.065 ;
      LAYER Metal2 ;
        RECT -2.870 -117.640 -2.490 -117.260 ;
        RECT -2.155 -120.715 -1.855 -113.675 ;
        RECT 0.870 -118.845 1.190 -113.685 ;
        RECT 6.880 -121.445 7.160 -118.410 ;
        RECT 9.630 -121.490 9.930 -114.335 ;
      LAYER Metal3 ;
        RECT -5.280 -117.575 -2.485 -117.280 ;
    END
  END b13_not
  PIN b13
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.270 -114.265 4.650 -113.885 ;
        RECT 2.670 -114.780 3.870 -114.490 ;
        RECT -2.860 -116.950 3.865 -116.650 ;
        RECT 3.460 -120.555 4.650 -120.270 ;
        RECT 2.680 -121.220 3.060 -120.840 ;
      LAYER Metal2 ;
        RECT -2.835 -116.970 -2.455 -116.590 ;
        RECT 2.720 -121.230 3.020 -114.420 ;
        RECT 3.510 -120.635 3.820 -114.445 ;
        RECT 4.305 -120.705 4.605 -113.875 ;
      LAYER Metal3 ;
        RECT -5.315 -116.945 -2.440 -116.650 ;
    END
  END b13
  PIN a13_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.590 -112.030 31.045 -111.650 ;
        RECT 29.750 -114.330 31.045 -113.950 ;
        RECT 43.235 -114.330 44.545 -113.950 ;
        RECT 28.080 -115.655 44.090 -115.280 ;
        RECT -2.880 -116.235 10.680 -115.935 ;
        RECT 12.585 -116.235 31.005 -115.935 ;
        RECT -0.415 -119.910 2.505 -119.610 ;
        RECT 6.050 -119.925 9.420 -119.625 ;
        RECT 15.045 -119.910 17.965 -119.610 ;
        RECT 21.510 -119.925 24.880 -119.625 ;
        RECT 29.760 -119.830 31.065 -119.450 ;
        RECT 43.100 -119.830 44.565 -119.450 ;
        RECT 29.575 -121.830 31.065 -121.450 ;
      LAYER Metal2 ;
        RECT -2.880 -116.285 -2.500 -115.905 ;
        RECT -0.380 -119.960 -0.080 -115.900 ;
        RECT 6.110 -119.975 6.390 -115.885 ;
        RECT 10.300 -116.285 10.680 -115.905 ;
        RECT 12.570 -116.285 12.950 -115.880 ;
        RECT 15.080 -119.960 15.380 -115.900 ;
        RECT 21.570 -119.975 21.850 -115.885 ;
        RECT 29.880 -121.885 30.235 -111.580 ;
        RECT 30.545 -116.280 30.890 -115.225 ;
        RECT 43.390 -120.110 43.720 -113.915 ;
      LAYER Metal3 ;
        RECT -5.320 -116.230 -2.475 -115.935 ;
        RECT 10.245 -116.255 12.985 -115.925 ;
    END
  END a13_not_f
  PIN a13_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.285 -111.930 54.565 -111.550 ;
        RECT 39.785 -114.330 40.970 -113.950 ;
        RECT 53.285 -114.330 54.300 -113.950 ;
        RECT -2.875 -115.490 10.690 -115.175 ;
        RECT 12.580 -115.490 26.405 -115.190 ;
        RECT 28.080 -117.010 54.310 -116.620 ;
        RECT -1.645 -118.145 2.485 -117.845 ;
        RECT 4.860 -118.195 9.360 -117.885 ;
        RECT 13.815 -118.145 17.945 -117.845 ;
        RECT 20.320 -118.195 24.820 -117.885 ;
        RECT 39.765 -119.830 41.125 -119.450 ;
        RECT 53.265 -119.830 54.445 -119.450 ;
        RECT 53.265 -121.830 54.340 -121.450 ;
      LAYER Metal2 ;
        RECT -2.870 -115.535 -2.490 -115.155 ;
        RECT 10.295 -115.535 10.675 -115.155 ;
        RECT 12.565 -115.535 12.945 -115.130 ;
        RECT 26.030 -115.535 26.390 -113.705 ;
        RECT 28.210 -117.055 28.625 -113.705 ;
        RECT 40.405 -113.965 40.715 -113.935 ;
        RECT 40.405 -120.065 40.720 -113.965 ;
        RECT 53.905 -122.060 54.235 -111.365 ;
      LAYER Metal3 ;
        RECT 25.975 -114.090 28.680 -113.750 ;
        RECT -5.280 -115.495 -2.455 -115.190 ;
        RECT 10.240 -115.505 12.985 -115.175 ;
    END
  END a13_f
  PIN b12_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -2.320 -94.305 1.055 -93.905 ;
        RECT 9.460 -94.955 9.840 -94.575 ;
        RECT -3.010 -97.810 1.115 -97.540 ;
        RECT 0.690 -98.985 7.080 -98.695 ;
        RECT -2.330 -100.900 -1.950 -100.520 ;
        RECT 6.670 -101.625 9.850 -101.305 ;
      LAYER Metal2 ;
        RECT -3.000 -97.880 -2.620 -97.500 ;
        RECT -2.285 -100.955 -1.985 -93.915 ;
        RECT 0.740 -99.085 1.060 -93.925 ;
        RECT 6.750 -101.685 7.030 -98.650 ;
        RECT 9.500 -101.730 9.800 -94.575 ;
      LAYER Metal3 ;
        RECT -5.410 -97.815 -2.615 -97.520 ;
    END
  END b12_not
  PIN b12
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.140 -94.505 4.520 -94.125 ;
        RECT 2.540 -95.020 3.740 -94.730 ;
        RECT -2.990 -97.190 3.735 -96.890 ;
        RECT 3.330 -100.795 4.520 -100.510 ;
        RECT 2.550 -101.460 2.930 -101.080 ;
      LAYER Metal2 ;
        RECT -2.965 -97.210 -2.585 -96.830 ;
        RECT 2.590 -101.470 2.890 -94.660 ;
        RECT 3.380 -100.875 3.690 -94.685 ;
        RECT 4.175 -100.945 4.475 -94.115 ;
      LAYER Metal3 ;
        RECT -5.445 -97.185 -2.570 -96.890 ;
    END
  END b12
  PIN a12_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.460 -92.270 30.915 -91.890 ;
        RECT 29.620 -94.570 30.915 -94.190 ;
        RECT 43.105 -94.570 44.415 -94.190 ;
        RECT 27.950 -95.895 43.960 -95.520 ;
        RECT -3.010 -96.475 10.550 -96.175 ;
        RECT 12.455 -96.475 30.875 -96.175 ;
        RECT -0.545 -100.150 2.375 -99.850 ;
        RECT 5.920 -100.165 9.290 -99.865 ;
        RECT 14.915 -100.150 17.835 -99.850 ;
        RECT 21.380 -100.165 24.750 -99.865 ;
        RECT 29.630 -100.070 30.935 -99.690 ;
        RECT 42.970 -100.070 44.435 -99.690 ;
        RECT 29.445 -102.070 30.935 -101.690 ;
      LAYER Metal2 ;
        RECT -3.010 -96.525 -2.630 -96.145 ;
        RECT -0.510 -100.200 -0.210 -96.140 ;
        RECT 5.980 -100.215 6.260 -96.125 ;
        RECT 10.170 -96.525 10.550 -96.145 ;
        RECT 12.440 -96.525 12.820 -96.120 ;
        RECT 14.950 -100.200 15.250 -96.140 ;
        RECT 21.440 -100.215 21.720 -96.125 ;
        RECT 29.750 -102.125 30.105 -91.820 ;
        RECT 30.415 -96.520 30.760 -95.465 ;
        RECT 43.260 -100.350 43.590 -94.155 ;
      LAYER Metal3 ;
        RECT -5.450 -96.470 -2.605 -96.175 ;
        RECT 10.115 -96.495 12.855 -96.165 ;
    END
  END a12_not_f
  PIN a12_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.155 -92.170 54.435 -91.790 ;
        RECT 39.655 -94.570 40.840 -94.190 ;
        RECT 53.155 -94.570 54.170 -94.190 ;
        RECT -3.005 -95.730 10.560 -95.415 ;
        RECT 12.450 -95.730 26.275 -95.430 ;
        RECT 27.950 -97.250 54.180 -96.860 ;
        RECT -1.775 -98.385 2.355 -98.085 ;
        RECT 4.730 -98.435 9.230 -98.125 ;
        RECT 13.685 -98.385 17.815 -98.085 ;
        RECT 20.190 -98.435 24.690 -98.125 ;
        RECT 39.635 -100.070 40.995 -99.690 ;
        RECT 53.135 -100.070 54.315 -99.690 ;
        RECT 53.135 -102.070 54.210 -101.690 ;
      LAYER Metal2 ;
        RECT -3.000 -95.775 -2.620 -95.395 ;
        RECT 10.165 -95.775 10.545 -95.395 ;
        RECT 12.435 -95.775 12.815 -95.370 ;
        RECT 25.900 -95.775 26.260 -93.945 ;
        RECT 28.080 -97.295 28.495 -93.945 ;
        RECT 40.275 -94.205 40.585 -94.175 ;
        RECT 40.275 -100.305 40.590 -94.205 ;
        RECT 53.775 -102.300 54.105 -91.605 ;
      LAYER Metal3 ;
        RECT 25.845 -94.330 28.550 -93.990 ;
        RECT -5.410 -95.735 -2.585 -95.430 ;
        RECT 10.110 -95.745 12.855 -95.415 ;
    END
  END a12_f
  PIN b11_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -2.190 -74.595 1.185 -74.195 ;
        RECT 9.590 -75.245 9.970 -74.865 ;
        RECT -2.880 -78.100 1.245 -77.830 ;
        RECT 0.820 -79.275 7.210 -78.985 ;
        RECT -2.200 -81.190 -1.820 -80.810 ;
        RECT 6.800 -81.915 9.980 -81.595 ;
      LAYER Metal2 ;
        RECT -2.870 -78.170 -2.490 -77.790 ;
        RECT -2.155 -81.245 -1.855 -74.205 ;
        RECT 0.870 -79.375 1.190 -74.215 ;
        RECT 6.880 -81.975 7.160 -78.940 ;
        RECT 9.630 -82.020 9.930 -74.865 ;
      LAYER Metal3 ;
        RECT -5.280 -78.105 -2.485 -77.810 ;
    END
  END b11_not
  PIN b11
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.270 -74.795 4.650 -74.415 ;
        RECT 2.670 -75.310 3.870 -75.020 ;
        RECT -2.860 -77.480 3.865 -77.180 ;
        RECT 3.460 -81.085 4.650 -80.800 ;
        RECT 2.680 -81.750 3.060 -81.370 ;
      LAYER Metal2 ;
        RECT -2.835 -77.500 -2.455 -77.120 ;
        RECT 2.720 -81.760 3.020 -74.950 ;
        RECT 3.510 -81.165 3.820 -74.975 ;
        RECT 4.305 -81.235 4.605 -74.405 ;
      LAYER Metal3 ;
        RECT -5.315 -77.475 -2.440 -77.180 ;
    END
  END b11
  PIN a11_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.590 -72.560 31.045 -72.180 ;
        RECT 29.750 -74.860 31.045 -74.480 ;
        RECT 43.235 -74.860 44.545 -74.480 ;
        RECT 28.080 -76.185 44.090 -75.810 ;
        RECT -2.880 -76.765 10.680 -76.465 ;
        RECT 12.585 -76.765 31.005 -76.465 ;
        RECT -0.415 -80.440 2.505 -80.140 ;
        RECT 6.050 -80.455 9.420 -80.155 ;
        RECT 15.045 -80.440 17.965 -80.140 ;
        RECT 21.510 -80.455 24.880 -80.155 ;
        RECT 29.760 -80.360 31.065 -79.980 ;
        RECT 43.100 -80.360 44.565 -79.980 ;
        RECT 29.575 -82.360 31.065 -81.980 ;
      LAYER Metal2 ;
        RECT -2.880 -76.815 -2.500 -76.435 ;
        RECT -0.380 -80.490 -0.080 -76.430 ;
        RECT 6.110 -80.505 6.390 -76.415 ;
        RECT 10.300 -76.815 10.680 -76.435 ;
        RECT 12.570 -76.815 12.950 -76.410 ;
        RECT 15.080 -80.490 15.380 -76.430 ;
        RECT 21.570 -80.505 21.850 -76.415 ;
        RECT 29.880 -82.415 30.235 -72.110 ;
        RECT 30.545 -76.810 30.890 -75.755 ;
        RECT 43.390 -80.640 43.720 -74.445 ;
      LAYER Metal3 ;
        RECT -5.320 -76.760 -2.475 -76.465 ;
        RECT 10.245 -76.785 12.985 -76.455 ;
    END
  END a11_not_f
  PIN a11_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.285 -72.460 54.565 -72.080 ;
        RECT 39.785 -74.860 40.970 -74.480 ;
        RECT 53.285 -74.860 54.300 -74.480 ;
        RECT -2.875 -76.020 10.690 -75.705 ;
        RECT 12.580 -76.020 26.405 -75.720 ;
        RECT 28.080 -77.540 54.310 -77.150 ;
        RECT -1.645 -78.675 2.485 -78.375 ;
        RECT 4.860 -78.725 9.360 -78.415 ;
        RECT 13.815 -78.675 17.945 -78.375 ;
        RECT 20.320 -78.725 24.820 -78.415 ;
        RECT 39.765 -80.360 41.125 -79.980 ;
        RECT 53.265 -80.360 54.445 -79.980 ;
        RECT 53.265 -82.360 54.340 -81.980 ;
      LAYER Metal2 ;
        RECT -2.870 -76.065 -2.490 -75.685 ;
        RECT 10.295 -76.065 10.675 -75.685 ;
        RECT 12.565 -76.065 12.945 -75.660 ;
        RECT 26.030 -76.065 26.390 -74.235 ;
        RECT 28.210 -77.585 28.625 -74.235 ;
        RECT 40.405 -74.495 40.715 -74.465 ;
        RECT 40.405 -80.595 40.720 -74.495 ;
        RECT 53.905 -82.590 54.235 -71.895 ;
      LAYER Metal3 ;
        RECT 25.975 -74.620 28.680 -74.280 ;
        RECT -5.280 -76.025 -2.455 -75.720 ;
        RECT 10.240 -76.035 12.985 -75.705 ;
    END
  END a11_f
  PIN b10_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -1.995 -54.755 1.380 -54.355 ;
        RECT 9.785 -55.405 10.165 -55.025 ;
        RECT -2.685 -58.260 1.440 -57.990 ;
        RECT 1.015 -59.435 7.405 -59.145 ;
        RECT -2.005 -61.350 -1.625 -60.970 ;
        RECT 6.995 -62.075 10.175 -61.755 ;
      LAYER Metal2 ;
        RECT -2.675 -58.330 -2.295 -57.950 ;
        RECT -1.960 -61.405 -1.660 -54.365 ;
        RECT 1.065 -59.535 1.385 -54.375 ;
        RECT 7.075 -62.135 7.355 -59.100 ;
        RECT 9.825 -62.180 10.125 -55.025 ;
      LAYER Metal3 ;
        RECT -5.085 -58.265 -2.290 -57.970 ;
    END
  END b10_not
  PIN b10
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.465 -54.955 4.845 -54.575 ;
        RECT 2.865 -55.470 4.065 -55.180 ;
        RECT -2.665 -57.640 4.060 -57.340 ;
        RECT 3.655 -61.245 4.845 -60.960 ;
        RECT 2.875 -61.910 3.255 -61.530 ;
      LAYER Metal2 ;
        RECT -2.640 -57.660 -2.260 -57.280 ;
        RECT 2.915 -61.920 3.215 -55.110 ;
        RECT 3.705 -61.325 4.015 -55.135 ;
        RECT 4.500 -61.395 4.800 -54.565 ;
      LAYER Metal3 ;
        RECT -5.120 -57.635 -2.245 -57.340 ;
    END
  END b10
  PIN a10_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.785 -52.720 31.240 -52.340 ;
        RECT 29.945 -55.020 31.240 -54.640 ;
        RECT 43.430 -55.020 44.740 -54.640 ;
        RECT 28.275 -56.345 44.285 -55.970 ;
        RECT -2.685 -56.925 10.875 -56.625 ;
        RECT 12.780 -56.925 31.200 -56.625 ;
        RECT -0.220 -60.600 2.700 -60.300 ;
        RECT 6.245 -60.615 9.615 -60.315 ;
        RECT 15.240 -60.600 18.160 -60.300 ;
        RECT 21.705 -60.615 25.075 -60.315 ;
        RECT 29.955 -60.520 31.260 -60.140 ;
        RECT 43.295 -60.520 44.760 -60.140 ;
        RECT 29.770 -62.520 31.260 -62.140 ;
      LAYER Metal2 ;
        RECT -2.685 -56.975 -2.305 -56.595 ;
        RECT -0.185 -60.650 0.115 -56.590 ;
        RECT 6.305 -60.665 6.585 -56.575 ;
        RECT 10.495 -56.975 10.875 -56.595 ;
        RECT 12.765 -56.975 13.145 -56.570 ;
        RECT 15.275 -60.650 15.575 -56.590 ;
        RECT 21.765 -60.665 22.045 -56.575 ;
        RECT 30.075 -62.575 30.430 -52.270 ;
        RECT 30.740 -56.970 31.085 -55.915 ;
        RECT 43.585 -60.800 43.915 -54.605 ;
      LAYER Metal3 ;
        RECT -5.125 -56.920 -2.280 -56.625 ;
        RECT 10.440 -56.945 13.180 -56.615 ;
    END
  END a10_not_f
  PIN a10_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.480 -52.620 54.760 -52.240 ;
        RECT 39.980 -55.020 41.165 -54.640 ;
        RECT 53.480 -55.020 54.495 -54.640 ;
        RECT -2.680 -56.180 10.885 -55.865 ;
        RECT 12.775 -56.180 26.600 -55.880 ;
        RECT 28.275 -57.700 54.505 -57.310 ;
        RECT -1.450 -58.835 2.680 -58.535 ;
        RECT 5.055 -58.885 9.555 -58.575 ;
        RECT 14.010 -58.835 18.140 -58.535 ;
        RECT 20.515 -58.885 25.015 -58.575 ;
        RECT 39.960 -60.520 41.320 -60.140 ;
        RECT 53.460 -60.520 54.640 -60.140 ;
        RECT 53.460 -62.520 54.535 -62.140 ;
      LAYER Metal2 ;
        RECT -2.675 -56.225 -2.295 -55.845 ;
        RECT 10.490 -56.225 10.870 -55.845 ;
        RECT 12.760 -56.225 13.140 -55.820 ;
        RECT 26.225 -56.225 26.585 -54.395 ;
        RECT 28.405 -57.745 28.820 -54.395 ;
        RECT 40.600 -54.655 40.910 -54.625 ;
        RECT 40.600 -60.755 40.915 -54.655 ;
        RECT 54.100 -62.750 54.430 -52.055 ;
      LAYER Metal3 ;
        RECT 26.170 -54.780 28.875 -54.440 ;
        RECT -5.085 -56.185 -2.260 -55.880 ;
        RECT 10.435 -56.195 13.180 -55.865 ;
    END
  END a10_f
  PIN b9_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -2.185 -35.045 1.190 -34.645 ;
        RECT 9.595 -35.695 9.975 -35.315 ;
        RECT -2.875 -38.550 1.250 -38.280 ;
        RECT 0.825 -39.725 7.215 -39.435 ;
        RECT -2.195 -41.640 -1.815 -41.260 ;
        RECT 6.805 -42.365 9.985 -42.045 ;
      LAYER Metal2 ;
        RECT -2.865 -38.620 -2.485 -38.240 ;
        RECT -2.150 -41.695 -1.850 -34.655 ;
        RECT 0.875 -39.825 1.195 -34.665 ;
        RECT 6.885 -42.425 7.165 -39.390 ;
        RECT 9.635 -42.470 9.935 -35.315 ;
      LAYER Metal3 ;
        RECT -5.275 -38.555 -2.480 -38.260 ;
    END
  END b9_not
  PIN b9
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.275 -35.245 4.655 -34.865 ;
        RECT 2.675 -35.760 3.875 -35.470 ;
        RECT -2.855 -37.930 3.870 -37.630 ;
        RECT 3.465 -41.535 4.655 -41.250 ;
        RECT 2.685 -42.200 3.065 -41.820 ;
      LAYER Metal2 ;
        RECT -2.830 -37.950 -2.450 -37.570 ;
        RECT 2.725 -42.210 3.025 -35.400 ;
        RECT 3.515 -41.615 3.825 -35.425 ;
        RECT 4.310 -41.685 4.610 -34.855 ;
      LAYER Metal3 ;
        RECT -5.310 -37.925 -2.435 -37.630 ;
    END
  END b9
  PIN a9_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.595 -33.010 31.050 -32.630 ;
        RECT 29.755 -35.310 31.050 -34.930 ;
        RECT 43.240 -35.310 44.550 -34.930 ;
        RECT 28.085 -36.635 44.095 -36.260 ;
        RECT -2.875 -37.215 10.685 -36.915 ;
        RECT 12.590 -37.215 31.010 -36.915 ;
        RECT -0.410 -40.890 2.510 -40.590 ;
        RECT 6.055 -40.905 9.425 -40.605 ;
        RECT 15.050 -40.890 17.970 -40.590 ;
        RECT 21.515 -40.905 24.885 -40.605 ;
        RECT 29.765 -40.810 31.070 -40.430 ;
        RECT 43.105 -40.810 44.570 -40.430 ;
        RECT 29.580 -42.810 31.070 -42.430 ;
      LAYER Metal2 ;
        RECT -2.875 -37.265 -2.495 -36.885 ;
        RECT -0.375 -40.940 -0.075 -36.880 ;
        RECT 6.115 -40.955 6.395 -36.865 ;
        RECT 10.305 -37.265 10.685 -36.885 ;
        RECT 12.575 -37.265 12.955 -36.860 ;
        RECT 15.085 -40.940 15.385 -36.880 ;
        RECT 21.575 -40.955 21.855 -36.865 ;
        RECT 29.885 -42.865 30.240 -32.560 ;
        RECT 30.550 -37.260 30.895 -36.205 ;
        RECT 43.395 -41.090 43.725 -34.895 ;
      LAYER Metal3 ;
        RECT -5.315 -37.210 -2.470 -36.915 ;
        RECT 10.250 -37.235 12.990 -36.905 ;
    END
  END a9_not_f
  PIN a9_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.290 -32.910 54.570 -32.530 ;
        RECT 39.790 -35.310 40.975 -34.930 ;
        RECT 53.290 -35.310 54.305 -34.930 ;
        RECT -2.870 -36.470 10.695 -36.155 ;
        RECT 12.585 -36.470 26.410 -36.170 ;
        RECT 28.085 -37.990 54.315 -37.600 ;
        RECT -1.640 -39.125 2.490 -38.825 ;
        RECT 4.865 -39.175 9.365 -38.865 ;
        RECT 13.820 -39.125 17.950 -38.825 ;
        RECT 20.325 -39.175 24.825 -38.865 ;
        RECT 39.770 -40.810 41.130 -40.430 ;
        RECT 53.270 -40.810 54.450 -40.430 ;
        RECT 53.270 -42.810 54.345 -42.430 ;
      LAYER Metal2 ;
        RECT -2.865 -36.515 -2.485 -36.135 ;
        RECT 10.300 -36.515 10.680 -36.135 ;
        RECT 12.570 -36.515 12.950 -36.110 ;
        RECT 26.035 -36.515 26.395 -34.685 ;
        RECT 28.215 -38.035 28.630 -34.685 ;
        RECT 40.410 -34.945 40.720 -34.915 ;
        RECT 40.410 -41.045 40.725 -34.945 ;
        RECT 53.910 -43.040 54.240 -32.345 ;
      LAYER Metal3 ;
        RECT 25.980 -35.070 28.685 -34.730 ;
        RECT -5.275 -36.475 -2.450 -36.170 ;
        RECT 10.245 -36.485 12.990 -36.155 ;
    END
  END a9_f
  PIN b8_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -2.140 -15.355 1.235 -14.955 ;
        RECT 9.640 -16.005 10.020 -15.625 ;
        RECT -2.830 -18.860 1.295 -18.590 ;
        RECT 0.870 -20.035 7.260 -19.745 ;
        RECT -2.150 -21.950 -1.770 -21.570 ;
        RECT 6.850 -22.675 10.030 -22.355 ;
      LAYER Metal2 ;
        RECT -2.820 -18.930 -2.440 -18.550 ;
        RECT -2.105 -22.005 -1.805 -14.965 ;
        RECT 0.920 -20.135 1.240 -14.975 ;
        RECT 6.930 -22.735 7.210 -19.700 ;
        RECT 9.680 -22.780 9.980 -15.625 ;
      LAYER Metal3 ;
        RECT -5.230 -18.865 -2.435 -18.570 ;
    END
  END b8_not
  PIN b8
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.320 -15.555 4.700 -15.175 ;
        RECT 2.720 -16.070 3.920 -15.780 ;
        RECT -2.810 -18.240 3.915 -17.940 ;
        RECT 3.510 -21.845 4.700 -21.560 ;
        RECT 2.730 -22.510 3.110 -22.130 ;
      LAYER Metal2 ;
        RECT -2.785 -18.260 -2.405 -17.880 ;
        RECT 2.770 -22.520 3.070 -15.710 ;
        RECT 3.560 -21.925 3.870 -15.735 ;
        RECT 4.355 -21.995 4.655 -15.165 ;
      LAYER Metal3 ;
        RECT -5.265 -18.235 -2.390 -17.940 ;
    END
  END b8
  PIN a8_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.640 -13.320 31.095 -12.940 ;
        RECT 29.800 -15.620 31.095 -15.240 ;
        RECT 43.285 -15.620 44.595 -15.240 ;
        RECT 28.130 -16.945 44.140 -16.570 ;
        RECT -2.830 -17.525 10.730 -17.225 ;
        RECT 12.635 -17.525 31.055 -17.225 ;
        RECT -0.365 -21.200 2.555 -20.900 ;
        RECT 6.100 -21.215 9.470 -20.915 ;
        RECT 15.095 -21.200 18.015 -20.900 ;
        RECT 21.560 -21.215 24.930 -20.915 ;
        RECT 29.810 -21.120 31.115 -20.740 ;
        RECT 43.150 -21.120 44.615 -20.740 ;
        RECT 29.625 -23.120 31.115 -22.740 ;
      LAYER Metal2 ;
        RECT -2.830 -17.575 -2.450 -17.195 ;
        RECT -0.330 -21.250 -0.030 -17.190 ;
        RECT 6.160 -21.265 6.440 -17.175 ;
        RECT 10.350 -17.575 10.730 -17.195 ;
        RECT 12.620 -17.575 13.000 -17.170 ;
        RECT 15.130 -21.250 15.430 -17.190 ;
        RECT 21.620 -21.265 21.900 -17.175 ;
        RECT 29.930 -23.175 30.285 -12.870 ;
        RECT 30.595 -17.570 30.940 -16.515 ;
        RECT 43.440 -21.400 43.770 -15.205 ;
      LAYER Metal3 ;
        RECT -5.270 -17.520 -2.425 -17.225 ;
        RECT 10.295 -17.545 13.035 -17.215 ;
    END
  END a8_not_f
  PIN a8_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.335 -13.220 54.615 -12.840 ;
        RECT 39.835 -15.620 41.020 -15.240 ;
        RECT 53.335 -15.620 54.350 -15.240 ;
        RECT -2.825 -16.780 10.740 -16.465 ;
        RECT 12.630 -16.780 26.455 -16.480 ;
        RECT 28.130 -18.300 54.360 -17.910 ;
        RECT -1.595 -19.435 2.535 -19.135 ;
        RECT 4.910 -19.485 9.410 -19.175 ;
        RECT 13.865 -19.435 17.995 -19.135 ;
        RECT 20.370 -19.485 24.870 -19.175 ;
        RECT 39.815 -21.120 41.175 -20.740 ;
        RECT 53.315 -21.120 54.495 -20.740 ;
        RECT 53.315 -23.120 54.390 -22.740 ;
      LAYER Metal2 ;
        RECT -2.820 -16.825 -2.440 -16.445 ;
        RECT 10.345 -16.825 10.725 -16.445 ;
        RECT 12.615 -16.825 12.995 -16.420 ;
        RECT 26.080 -16.825 26.440 -14.995 ;
        RECT 28.260 -18.345 28.675 -14.995 ;
        RECT 40.455 -15.255 40.765 -15.225 ;
        RECT 40.455 -21.355 40.770 -15.255 ;
        RECT 53.955 -23.350 54.285 -12.655 ;
      LAYER Metal3 ;
        RECT 26.025 -15.380 28.730 -15.040 ;
        RECT -5.230 -16.785 -2.405 -16.480 ;
        RECT 10.290 -16.795 13.035 -16.465 ;
    END
  END a8_f
  PIN b7_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -2.290 4.440 1.085 4.840 ;
        RECT 9.490 3.790 9.870 4.170 ;
        RECT -2.980 0.935 1.145 1.205 ;
        RECT 0.720 -0.240 7.110 0.050 ;
        RECT -2.300 -2.155 -1.920 -1.775 ;
        RECT 6.700 -2.880 9.880 -2.560 ;
      LAYER Metal2 ;
        RECT -2.970 0.865 -2.590 1.245 ;
        RECT -2.255 -2.210 -1.955 4.830 ;
        RECT 0.770 -0.340 1.090 4.820 ;
        RECT 6.780 -2.940 7.060 0.095 ;
        RECT 9.530 -2.985 9.830 4.170 ;
      LAYER Metal3 ;
        RECT -5.380 0.930 -2.585 1.225 ;
    END
  END b7_not
  PIN b7
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.170 4.240 4.550 4.620 ;
        RECT 2.570 3.725 3.770 4.015 ;
        RECT -2.960 1.555 3.765 1.855 ;
        RECT 3.360 -2.050 4.550 -1.765 ;
        RECT 2.580 -2.715 2.960 -2.335 ;
      LAYER Metal2 ;
        RECT -2.935 1.535 -2.555 1.915 ;
        RECT 2.620 -2.725 2.920 4.085 ;
        RECT 3.410 -2.130 3.720 4.060 ;
        RECT 4.205 -2.200 4.505 4.630 ;
      LAYER Metal3 ;
        RECT -5.415 1.560 -2.540 1.855 ;
    END
  END b7
  PIN a7_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.490 6.475 30.945 6.855 ;
        RECT 29.650 4.175 30.945 4.555 ;
        RECT 43.135 4.175 44.445 4.555 ;
        RECT 27.980 2.850 43.990 3.225 ;
        RECT -2.980 2.270 10.580 2.570 ;
        RECT 12.485 2.270 30.905 2.570 ;
        RECT -0.515 -1.405 2.405 -1.105 ;
        RECT 5.950 -1.420 9.320 -1.120 ;
        RECT 14.945 -1.405 17.865 -1.105 ;
        RECT 21.410 -1.420 24.780 -1.120 ;
        RECT 29.660 -1.325 30.965 -0.945 ;
        RECT 43.000 -1.325 44.465 -0.945 ;
        RECT 29.475 -3.325 30.965 -2.945 ;
      LAYER Metal2 ;
        RECT -2.980 2.220 -2.600 2.600 ;
        RECT -0.480 -1.455 -0.180 2.605 ;
        RECT 6.010 -1.470 6.290 2.620 ;
        RECT 10.200 2.220 10.580 2.600 ;
        RECT 12.470 2.220 12.850 2.625 ;
        RECT 14.980 -1.455 15.280 2.605 ;
        RECT 21.470 -1.470 21.750 2.620 ;
        RECT 29.780 -3.380 30.135 6.925 ;
        RECT 30.445 2.225 30.790 3.280 ;
        RECT 43.290 -1.605 43.620 4.590 ;
      LAYER Metal3 ;
        RECT -5.420 2.275 -2.575 2.570 ;
        RECT 10.145 2.250 12.885 2.580 ;
    END
  END a7_not_f
  PIN a7_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.185 6.575 54.465 6.955 ;
        RECT 39.685 4.175 40.870 4.555 ;
        RECT 53.185 4.175 54.200 4.555 ;
        RECT -2.975 3.015 10.590 3.330 ;
        RECT 12.480 3.015 26.305 3.315 ;
        RECT 27.980 1.495 54.210 1.885 ;
        RECT -1.745 0.360 2.385 0.660 ;
        RECT 4.760 0.310 9.260 0.620 ;
        RECT 13.715 0.360 17.845 0.660 ;
        RECT 20.220 0.310 24.720 0.620 ;
        RECT 39.665 -1.325 41.025 -0.945 ;
        RECT 53.165 -1.325 54.345 -0.945 ;
        RECT 53.165 -3.325 54.240 -2.945 ;
      LAYER Metal2 ;
        RECT -2.970 2.970 -2.590 3.350 ;
        RECT 10.195 2.970 10.575 3.350 ;
        RECT 12.465 2.970 12.845 3.375 ;
        RECT 25.930 2.970 26.290 4.800 ;
        RECT 28.110 1.450 28.525 4.800 ;
        RECT 40.305 4.540 40.615 4.570 ;
        RECT 40.305 -1.560 40.620 4.540 ;
        RECT 53.805 -3.555 54.135 7.140 ;
      LAYER Metal3 ;
        RECT 25.875 4.415 28.580 4.755 ;
        RECT -5.380 3.010 -2.555 3.315 ;
        RECT 10.140 3.000 12.885 3.330 ;
    END
  END a7_f
  PIN b6_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -2.260 24.235 1.115 24.635 ;
        RECT 9.520 23.585 9.900 23.965 ;
        RECT -2.950 20.730 1.175 21.000 ;
        RECT 0.750 19.555 7.140 19.845 ;
        RECT -2.270 17.640 -1.890 18.020 ;
        RECT 6.730 16.915 9.910 17.235 ;
      LAYER Metal2 ;
        RECT -2.940 20.660 -2.560 21.040 ;
        RECT -2.225 17.585 -1.925 24.625 ;
        RECT 0.800 19.455 1.120 24.615 ;
        RECT 6.810 16.855 7.090 19.890 ;
        RECT 9.560 16.810 9.860 23.965 ;
      LAYER Metal3 ;
        RECT -5.350 20.725 -2.555 21.020 ;
    END
  END b6_not
  PIN b6
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.200 24.035 4.580 24.415 ;
        RECT 2.600 23.520 3.800 23.810 ;
        RECT -2.930 21.350 3.795 21.650 ;
        RECT 3.390 17.745 4.580 18.030 ;
        RECT 2.610 17.080 2.990 17.460 ;
      LAYER Metal2 ;
        RECT -2.905 21.330 -2.525 21.710 ;
        RECT 2.650 17.070 2.950 23.880 ;
        RECT 3.440 17.665 3.750 23.855 ;
        RECT 4.235 17.595 4.535 24.425 ;
      LAYER Metal3 ;
        RECT -5.385 21.355 -2.510 21.650 ;
    END
  END b6
  PIN a6_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.520 26.270 30.975 26.650 ;
        RECT 29.680 23.970 30.975 24.350 ;
        RECT 43.165 23.970 44.475 24.350 ;
        RECT 28.010 22.645 44.020 23.020 ;
        RECT -2.950 22.065 10.610 22.365 ;
        RECT 12.515 22.065 30.935 22.365 ;
        RECT -0.485 18.390 2.435 18.690 ;
        RECT 5.980 18.375 9.350 18.675 ;
        RECT 14.975 18.390 17.895 18.690 ;
        RECT 21.440 18.375 24.810 18.675 ;
        RECT 29.690 18.470 30.995 18.850 ;
        RECT 43.030 18.470 44.495 18.850 ;
        RECT 29.505 16.470 30.995 16.850 ;
      LAYER Metal2 ;
        RECT -2.950 22.015 -2.570 22.395 ;
        RECT -0.450 18.340 -0.150 22.400 ;
        RECT 6.040 18.325 6.320 22.415 ;
        RECT 10.230 22.015 10.610 22.395 ;
        RECT 12.500 22.015 12.880 22.420 ;
        RECT 15.010 18.340 15.310 22.400 ;
        RECT 21.500 18.325 21.780 22.415 ;
        RECT 29.810 16.415 30.165 26.720 ;
        RECT 30.475 22.020 30.820 23.075 ;
        RECT 43.320 18.190 43.650 24.385 ;
      LAYER Metal3 ;
        RECT -5.390 22.070 -2.545 22.365 ;
        RECT 10.175 22.045 12.915 22.375 ;
    END
  END a6_not_f
  PIN a6_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.215 26.370 54.495 26.750 ;
        RECT 39.715 23.970 40.900 24.350 ;
        RECT 53.215 23.970 54.230 24.350 ;
        RECT -2.945 22.810 10.620 23.125 ;
        RECT 12.510 22.810 26.335 23.110 ;
        RECT 28.010 21.290 54.240 21.680 ;
        RECT -1.715 20.155 2.415 20.455 ;
        RECT 4.790 20.105 9.290 20.415 ;
        RECT 13.745 20.155 17.875 20.455 ;
        RECT 20.250 20.105 24.750 20.415 ;
        RECT 39.695 18.470 41.055 18.850 ;
        RECT 53.195 18.470 54.375 18.850 ;
        RECT 53.195 16.470 54.270 16.850 ;
      LAYER Metal2 ;
        RECT -2.940 22.765 -2.560 23.145 ;
        RECT 10.225 22.765 10.605 23.145 ;
        RECT 12.495 22.765 12.875 23.170 ;
        RECT 25.960 22.765 26.320 24.595 ;
        RECT 28.140 21.245 28.555 24.595 ;
        RECT 40.335 24.335 40.645 24.365 ;
        RECT 40.335 18.235 40.650 24.335 ;
        RECT 53.835 16.240 54.165 26.935 ;
      LAYER Metal3 ;
        RECT 25.905 24.210 28.610 24.550 ;
        RECT -5.350 22.805 -2.525 23.110 ;
        RECT 10.170 22.795 12.915 23.125 ;
    END
  END a6_f
  PIN b5_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -2.210 44.045 1.165 44.445 ;
        RECT 9.570 43.395 9.950 43.775 ;
        RECT -2.900 40.540 1.225 40.810 ;
        RECT 0.800 39.365 7.190 39.655 ;
        RECT -2.220 37.450 -1.840 37.830 ;
        RECT 6.780 36.725 9.960 37.045 ;
      LAYER Metal2 ;
        RECT -2.890 40.470 -2.510 40.850 ;
        RECT -2.175 37.395 -1.875 44.435 ;
        RECT 0.850 39.265 1.170 44.425 ;
        RECT 6.860 36.665 7.140 39.700 ;
        RECT 9.610 36.620 9.910 43.775 ;
      LAYER Metal3 ;
        RECT -5.300 40.535 -2.505 40.830 ;
    END
  END b5_not
  PIN b5
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.250 43.845 4.630 44.225 ;
        RECT 2.650 43.330 3.850 43.620 ;
        RECT -2.880 41.160 3.845 41.460 ;
        RECT 3.440 37.555 4.630 37.840 ;
        RECT 2.660 36.890 3.040 37.270 ;
      LAYER Metal2 ;
        RECT -2.855 41.140 -2.475 41.520 ;
        RECT 2.700 36.880 3.000 43.690 ;
        RECT 3.490 37.475 3.800 43.665 ;
        RECT 4.285 37.405 4.585 44.235 ;
      LAYER Metal3 ;
        RECT -5.335 41.165 -2.460 41.460 ;
    END
  END b5
  PIN a5_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.570 46.080 31.025 46.460 ;
        RECT 29.730 43.780 31.025 44.160 ;
        RECT 43.215 43.780 44.525 44.160 ;
        RECT 28.060 42.455 44.070 42.830 ;
        RECT -2.900 41.875 10.660 42.175 ;
        RECT 12.565 41.875 30.985 42.175 ;
        RECT -0.435 38.200 2.485 38.500 ;
        RECT 6.030 38.185 9.400 38.485 ;
        RECT 15.025 38.200 17.945 38.500 ;
        RECT 21.490 38.185 24.860 38.485 ;
        RECT 29.740 38.280 31.045 38.660 ;
        RECT 43.080 38.280 44.545 38.660 ;
        RECT 29.555 36.280 31.045 36.660 ;
      LAYER Metal2 ;
        RECT -2.900 41.825 -2.520 42.205 ;
        RECT -0.400 38.150 -0.100 42.210 ;
        RECT 6.090 38.135 6.370 42.225 ;
        RECT 10.280 41.825 10.660 42.205 ;
        RECT 12.550 41.825 12.930 42.230 ;
        RECT 15.060 38.150 15.360 42.210 ;
        RECT 21.550 38.135 21.830 42.225 ;
        RECT 29.860 36.225 30.215 46.530 ;
        RECT 30.525 41.830 30.870 42.885 ;
        RECT 43.370 38.000 43.700 44.195 ;
      LAYER Metal3 ;
        RECT -5.340 41.880 -2.495 42.175 ;
        RECT 10.225 41.855 12.965 42.185 ;
    END
  END a5_not_f
  PIN a5_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.265 46.180 54.545 46.560 ;
        RECT 39.765 43.780 40.950 44.160 ;
        RECT 53.265 43.780 54.280 44.160 ;
        RECT -2.895 42.620 10.670 42.935 ;
        RECT 12.560 42.620 26.385 42.920 ;
        RECT 28.060 41.100 54.290 41.490 ;
        RECT -1.665 39.965 2.465 40.265 ;
        RECT 4.840 39.915 9.340 40.225 ;
        RECT 13.795 39.965 17.925 40.265 ;
        RECT 20.300 39.915 24.800 40.225 ;
        RECT 39.745 38.280 41.105 38.660 ;
        RECT 53.245 38.280 54.425 38.660 ;
        RECT 53.245 36.280 54.320 36.660 ;
      LAYER Metal2 ;
        RECT -2.890 42.575 -2.510 42.955 ;
        RECT 10.275 42.575 10.655 42.955 ;
        RECT 12.545 42.575 12.925 42.980 ;
        RECT 26.010 42.575 26.370 44.405 ;
        RECT 28.190 41.055 28.605 44.405 ;
        RECT 40.385 44.145 40.695 44.175 ;
        RECT 40.385 38.045 40.700 44.145 ;
        RECT 53.885 36.050 54.215 46.745 ;
      LAYER Metal3 ;
        RECT 25.955 44.020 28.660 44.360 ;
        RECT -5.300 42.615 -2.475 42.920 ;
        RECT 10.220 42.605 12.965 42.935 ;
    END
  END a5_f
  PIN b4_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -2.340 63.805 1.035 64.205 ;
        RECT 9.440 63.155 9.820 63.535 ;
        RECT -3.030 60.300 1.095 60.570 ;
        RECT 0.670 59.125 7.060 59.415 ;
        RECT -2.350 57.210 -1.970 57.590 ;
        RECT 6.650 56.485 9.830 56.805 ;
      LAYER Metal2 ;
        RECT -3.020 60.230 -2.640 60.610 ;
        RECT -2.305 57.155 -2.005 64.195 ;
        RECT 0.720 59.025 1.040 64.185 ;
        RECT 6.730 56.425 7.010 59.460 ;
        RECT 9.480 56.380 9.780 63.535 ;
      LAYER Metal3 ;
        RECT -5.430 60.295 -2.635 60.590 ;
    END
  END b4_not
  PIN b4
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.120 63.605 4.500 63.985 ;
        RECT 2.520 63.090 3.720 63.380 ;
        RECT -3.010 60.920 3.715 61.220 ;
        RECT 3.310 57.315 4.500 57.600 ;
        RECT 2.530 56.650 2.910 57.030 ;
      LAYER Metal2 ;
        RECT -2.985 60.900 -2.605 61.280 ;
        RECT 2.570 56.640 2.870 63.450 ;
        RECT 3.360 57.235 3.670 63.425 ;
        RECT 4.155 57.165 4.455 63.995 ;
      LAYER Metal3 ;
        RECT -5.465 60.925 -2.590 61.220 ;
    END
  END b4
  PIN a4_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.440 65.840 30.895 66.220 ;
        RECT 29.600 63.540 30.895 63.920 ;
        RECT 43.085 63.540 44.395 63.920 ;
        RECT 27.930 62.215 43.940 62.590 ;
        RECT -3.030 61.635 10.530 61.935 ;
        RECT 12.435 61.635 30.855 61.935 ;
        RECT -0.565 57.960 2.355 58.260 ;
        RECT 5.900 57.945 9.270 58.245 ;
        RECT 14.895 57.960 17.815 58.260 ;
        RECT 21.360 57.945 24.730 58.245 ;
        RECT 29.610 58.040 30.915 58.420 ;
        RECT 42.950 58.040 44.415 58.420 ;
        RECT 29.425 56.040 30.915 56.420 ;
      LAYER Metal2 ;
        RECT -3.030 61.585 -2.650 61.965 ;
        RECT -0.530 57.910 -0.230 61.970 ;
        RECT 5.960 57.895 6.240 61.985 ;
        RECT 10.150 61.585 10.530 61.965 ;
        RECT 12.420 61.585 12.800 61.990 ;
        RECT 14.930 57.910 15.230 61.970 ;
        RECT 21.420 57.895 21.700 61.985 ;
        RECT 29.730 55.985 30.085 66.290 ;
        RECT 30.395 61.590 30.740 62.645 ;
        RECT 43.240 57.760 43.570 63.955 ;
      LAYER Metal3 ;
        RECT -5.470 61.640 -2.625 61.935 ;
        RECT 10.095 61.615 12.835 61.945 ;
    END
  END a4_not_f
  PIN a4_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.135 65.940 54.415 66.320 ;
        RECT 39.635 63.540 40.820 63.920 ;
        RECT 53.135 63.540 54.150 63.920 ;
        RECT -3.025 62.380 10.540 62.695 ;
        RECT 12.430 62.380 26.255 62.680 ;
        RECT 27.930 60.860 54.160 61.250 ;
        RECT -1.795 59.725 2.335 60.025 ;
        RECT 4.710 59.675 9.210 59.985 ;
        RECT 13.665 59.725 17.795 60.025 ;
        RECT 20.170 59.675 24.670 59.985 ;
        RECT 39.615 58.040 40.975 58.420 ;
        RECT 53.115 58.040 54.295 58.420 ;
        RECT 53.115 56.040 54.190 56.420 ;
      LAYER Metal2 ;
        RECT -3.020 62.335 -2.640 62.715 ;
        RECT 10.145 62.335 10.525 62.715 ;
        RECT 12.415 62.335 12.795 62.740 ;
        RECT 25.880 62.335 26.240 64.165 ;
        RECT 28.060 60.815 28.475 64.165 ;
        RECT 40.255 63.905 40.565 63.935 ;
        RECT 40.255 57.805 40.570 63.905 ;
        RECT 53.755 55.810 54.085 66.505 ;
      LAYER Metal3 ;
        RECT 25.825 63.780 28.530 64.120 ;
        RECT -5.430 62.375 -2.605 62.680 ;
        RECT 10.090 62.365 12.835 62.695 ;
    END
  END a4_f
  PIN b3_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -2.210 83.515 1.165 83.915 ;
        RECT 9.570 82.865 9.950 83.245 ;
        RECT -2.900 80.010 1.225 80.280 ;
        RECT 0.800 78.835 7.190 79.125 ;
        RECT -2.220 76.920 -1.840 77.300 ;
        RECT 6.780 76.195 9.960 76.515 ;
      LAYER Metal2 ;
        RECT -2.890 79.940 -2.510 80.320 ;
        RECT -2.175 76.865 -1.875 83.905 ;
        RECT 0.850 78.735 1.170 83.895 ;
        RECT 6.860 76.135 7.140 79.170 ;
        RECT 9.610 76.090 9.910 83.245 ;
      LAYER Metal3 ;
        RECT -5.300 80.005 -2.505 80.300 ;
    END
  END b3_not
  PIN b3
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.250 83.315 4.630 83.695 ;
        RECT 2.650 82.800 3.850 83.090 ;
        RECT -2.880 80.630 3.845 80.930 ;
        RECT 3.440 77.025 4.630 77.310 ;
        RECT 2.660 76.360 3.040 76.740 ;
      LAYER Metal2 ;
        RECT -2.855 80.610 -2.475 80.990 ;
        RECT 2.700 76.350 3.000 83.160 ;
        RECT 3.490 76.945 3.800 83.135 ;
        RECT 4.285 76.875 4.585 83.705 ;
      LAYER Metal3 ;
        RECT -5.335 80.635 -2.460 80.930 ;
    END
  END b3
  PIN a3_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.570 85.550 31.025 85.930 ;
        RECT 29.730 83.250 31.025 83.630 ;
        RECT 43.215 83.250 44.525 83.630 ;
        RECT 28.060 81.925 44.070 82.300 ;
        RECT -2.900 81.345 10.660 81.645 ;
        RECT 12.565 81.345 30.985 81.645 ;
        RECT -0.435 77.670 2.485 77.970 ;
        RECT 6.030 77.655 9.400 77.955 ;
        RECT 15.025 77.670 17.945 77.970 ;
        RECT 21.490 77.655 24.860 77.955 ;
        RECT 29.740 77.750 31.045 78.130 ;
        RECT 43.080 77.750 44.545 78.130 ;
        RECT 29.555 75.750 31.045 76.130 ;
      LAYER Metal2 ;
        RECT -2.900 81.295 -2.520 81.675 ;
        RECT -0.400 77.620 -0.100 81.680 ;
        RECT 6.090 77.605 6.370 81.695 ;
        RECT 10.280 81.295 10.660 81.675 ;
        RECT 12.550 81.295 12.930 81.700 ;
        RECT 15.060 77.620 15.360 81.680 ;
        RECT 21.550 77.605 21.830 81.695 ;
        RECT 29.860 75.695 30.215 86.000 ;
        RECT 30.525 81.300 30.870 82.355 ;
        RECT 43.370 77.470 43.700 83.665 ;
      LAYER Metal3 ;
        RECT -5.340 81.350 -2.495 81.645 ;
        RECT 10.225 81.325 12.965 81.655 ;
    END
  END a3_not_f
  PIN a3_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.265 85.650 54.545 86.030 ;
        RECT 39.765 83.250 40.950 83.630 ;
        RECT 53.265 83.250 54.280 83.630 ;
        RECT -2.895 82.090 10.670 82.405 ;
        RECT 12.560 82.090 26.385 82.390 ;
        RECT 28.060 80.570 54.290 80.960 ;
        RECT -1.665 79.435 2.465 79.735 ;
        RECT 4.840 79.385 9.340 79.695 ;
        RECT 13.795 79.435 17.925 79.735 ;
        RECT 20.300 79.385 24.800 79.695 ;
        RECT 39.745 77.750 41.105 78.130 ;
        RECT 53.245 77.750 54.425 78.130 ;
        RECT 53.245 75.750 54.320 76.130 ;
      LAYER Metal2 ;
        RECT -2.890 82.045 -2.510 82.425 ;
        RECT 10.275 82.045 10.655 82.425 ;
        RECT 12.545 82.045 12.925 82.450 ;
        RECT 26.010 82.045 26.370 83.875 ;
        RECT 28.190 80.525 28.605 83.875 ;
        RECT 40.385 83.615 40.695 83.645 ;
        RECT 40.385 77.515 40.700 83.615 ;
        RECT 53.885 75.520 54.215 86.215 ;
      LAYER Metal3 ;
        RECT 25.955 83.490 28.660 83.830 ;
        RECT -5.300 82.085 -2.475 82.390 ;
        RECT 10.220 82.075 12.965 82.405 ;
    END
  END a3_f
  PIN a0_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.315 144.890 54.595 145.270 ;
        RECT 39.815 142.490 41.000 142.870 ;
        RECT 53.315 142.490 54.330 142.870 ;
        RECT -2.845 141.330 10.720 141.645 ;
        RECT 12.610 141.330 26.435 141.630 ;
        RECT 28.110 139.810 54.340 140.200 ;
        RECT -1.615 138.675 2.515 138.975 ;
        RECT 4.890 138.625 9.390 138.935 ;
        RECT 13.845 138.675 17.975 138.975 ;
        RECT 20.350 138.625 24.850 138.935 ;
        RECT 39.795 136.990 41.155 137.370 ;
        RECT 53.295 136.990 54.475 137.370 ;
        RECT 53.295 134.990 54.370 135.370 ;
      LAYER Metal2 ;
        RECT -2.840 141.285 -2.460 141.665 ;
        RECT 10.325 141.285 10.705 141.665 ;
        RECT 12.595 141.285 12.975 141.690 ;
        RECT 26.060 141.285 26.420 143.115 ;
        RECT 28.240 139.765 28.655 143.115 ;
        RECT 40.435 142.855 40.745 142.885 ;
        RECT 40.435 136.755 40.750 142.855 ;
        RECT 53.935 134.760 54.265 145.455 ;
      LAYER Metal3 ;
        RECT 26.005 142.730 28.710 143.070 ;
        RECT -5.250 141.325 -2.425 141.630 ;
        RECT 10.270 141.315 13.015 141.645 ;
    END
  END a0_f
  PIN a0_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.620 144.790 31.075 145.170 ;
        RECT 29.780 142.490 31.075 142.870 ;
        RECT 43.265 142.490 44.575 142.870 ;
        RECT 28.110 141.165 44.120 141.540 ;
        RECT -2.850 140.585 10.710 140.885 ;
        RECT 12.615 140.585 31.035 140.885 ;
        RECT -0.385 136.910 2.535 137.210 ;
        RECT 6.080 136.895 9.450 137.195 ;
        RECT 15.075 136.910 17.995 137.210 ;
        RECT 21.540 136.895 24.910 137.195 ;
        RECT 29.790 136.990 31.095 137.370 ;
        RECT 43.130 136.990 44.595 137.370 ;
        RECT 29.605 134.990 31.095 135.370 ;
      LAYER Metal2 ;
        RECT -2.850 140.535 -2.470 140.915 ;
        RECT -0.350 136.860 -0.050 140.920 ;
        RECT 6.140 136.845 6.420 140.935 ;
        RECT 10.330 140.535 10.710 140.915 ;
        RECT 12.600 140.535 12.980 140.940 ;
        RECT 15.110 136.860 15.410 140.920 ;
        RECT 21.600 136.845 21.880 140.935 ;
        RECT 29.910 134.935 30.265 145.240 ;
        RECT 30.575 140.540 30.920 141.595 ;
        RECT 43.420 136.710 43.750 142.905 ;
      LAYER Metal3 ;
        RECT -5.290 140.590 -2.445 140.885 ;
        RECT 10.275 140.565 13.015 140.895 ;
    END
  END a0_not_f
  PIN b0
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.300 142.555 4.680 142.935 ;
        RECT 2.700 142.040 3.900 142.330 ;
        RECT -2.830 139.870 3.895 140.170 ;
        RECT 3.490 136.265 4.680 136.550 ;
        RECT 2.710 135.600 3.090 135.980 ;
      LAYER Metal2 ;
        RECT -2.805 139.850 -2.425 140.230 ;
        RECT 2.750 135.590 3.050 142.400 ;
        RECT 3.540 136.185 3.850 142.375 ;
        RECT 4.335 136.115 4.635 142.945 ;
      LAYER Metal3 ;
        RECT -5.285 139.875 -2.410 140.170 ;
    END
  END b0
  PIN b0_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -2.160 142.755 1.215 143.155 ;
        RECT 9.620 142.105 10.000 142.485 ;
        RECT -2.850 139.250 1.275 139.520 ;
        RECT 0.850 138.075 7.240 138.365 ;
        RECT -2.170 136.160 -1.790 136.540 ;
        RECT 6.830 135.435 10.010 135.755 ;
      LAYER Metal2 ;
        RECT -2.840 139.180 -2.460 139.560 ;
        RECT -2.125 136.105 -1.825 143.145 ;
        RECT 0.900 137.975 1.220 143.135 ;
        RECT 6.910 135.375 7.190 138.410 ;
        RECT 9.660 135.330 9.960 142.485 ;
      LAYER Metal3 ;
        RECT -5.250 139.245 -2.455 139.540 ;
    END
  END b0_not
  PIN b2_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -2.015 103.355 1.360 103.755 ;
        RECT 9.765 102.705 10.145 103.085 ;
        RECT -2.705 99.850 1.420 100.120 ;
        RECT 0.995 98.675 7.385 98.965 ;
        RECT -2.025 96.760 -1.645 97.140 ;
        RECT 6.975 96.035 10.155 96.355 ;
      LAYER Metal2 ;
        RECT -2.695 99.780 -2.315 100.160 ;
        RECT -1.980 96.705 -1.680 103.745 ;
        RECT 1.045 98.575 1.365 103.735 ;
        RECT 7.055 95.975 7.335 99.010 ;
        RECT 9.805 95.930 10.105 103.085 ;
      LAYER Metal3 ;
        RECT -5.105 99.845 -2.310 100.140 ;
    END
  END b2_not
  PIN b2
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.445 103.155 4.825 103.535 ;
        RECT 2.845 102.640 4.045 102.930 ;
        RECT -2.685 100.470 4.040 100.770 ;
        RECT 3.635 96.865 4.825 97.150 ;
        RECT 2.855 96.200 3.235 96.580 ;
      LAYER Metal2 ;
        RECT -2.660 100.450 -2.280 100.830 ;
        RECT 2.895 96.190 3.195 103.000 ;
        RECT 3.685 96.785 3.995 102.975 ;
        RECT 4.480 96.715 4.780 103.545 ;
      LAYER Metal3 ;
        RECT -5.140 100.475 -2.265 100.770 ;
    END
  END b2
  PIN a2_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.765 105.390 31.220 105.770 ;
        RECT 29.925 103.090 31.220 103.470 ;
        RECT 43.410 103.090 44.720 103.470 ;
        RECT 28.255 101.765 44.265 102.140 ;
        RECT -2.705 101.185 10.855 101.485 ;
        RECT 12.760 101.185 31.180 101.485 ;
        RECT -0.240 97.510 2.680 97.810 ;
        RECT 6.225 97.495 9.595 97.795 ;
        RECT 15.220 97.510 18.140 97.810 ;
        RECT 21.685 97.495 25.055 97.795 ;
        RECT 29.935 97.590 31.240 97.970 ;
        RECT 43.275 97.590 44.740 97.970 ;
        RECT 29.750 95.590 31.240 95.970 ;
      LAYER Metal2 ;
        RECT -2.705 101.135 -2.325 101.515 ;
        RECT -0.205 97.460 0.095 101.520 ;
        RECT 6.285 97.445 6.565 101.535 ;
        RECT 10.475 101.135 10.855 101.515 ;
        RECT 12.745 101.135 13.125 101.540 ;
        RECT 15.255 97.460 15.555 101.520 ;
        RECT 21.745 97.445 22.025 101.535 ;
        RECT 30.055 95.535 30.410 105.840 ;
        RECT 30.720 101.140 31.065 102.195 ;
        RECT 43.565 97.310 43.895 103.505 ;
      LAYER Metal3 ;
        RECT -5.145 101.190 -2.300 101.485 ;
        RECT 10.420 101.165 13.160 101.495 ;
    END
  END a2_not_f
  PIN a2_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.460 105.490 54.740 105.870 ;
        RECT 39.960 103.090 41.145 103.470 ;
        RECT 53.460 103.090 54.475 103.470 ;
        RECT -2.700 101.930 10.865 102.245 ;
        RECT 12.755 101.930 26.580 102.230 ;
        RECT 28.255 100.410 54.485 100.800 ;
        RECT -1.470 99.275 2.660 99.575 ;
        RECT 5.035 99.225 9.535 99.535 ;
        RECT 13.990 99.275 18.120 99.575 ;
        RECT 20.495 99.225 24.995 99.535 ;
        RECT 39.940 97.590 41.300 97.970 ;
        RECT 53.440 97.590 54.620 97.970 ;
        RECT 53.440 95.590 54.515 95.970 ;
      LAYER Metal2 ;
        RECT -2.695 101.885 -2.315 102.265 ;
        RECT 10.470 101.885 10.850 102.265 ;
        RECT 12.740 101.885 13.120 102.290 ;
        RECT 26.205 101.885 26.565 103.715 ;
        RECT 28.385 100.365 28.800 103.715 ;
        RECT 40.580 103.455 40.890 103.485 ;
        RECT 40.580 97.355 40.895 103.455 ;
        RECT 54.080 95.360 54.410 106.055 ;
      LAYER Metal3 ;
        RECT 26.150 103.330 28.855 103.670 ;
        RECT -5.105 101.925 -2.280 102.230 ;
        RECT 10.415 101.915 13.160 102.245 ;
    END
  END a2_f
  PIN b1_not
    ANTENNADIFFAREA 2.638650 ;
    PORT
      LAYER Metal1 ;
        RECT -2.205 123.065 1.170 123.465 ;
        RECT 9.575 122.415 9.955 122.795 ;
        RECT -2.895 119.560 1.230 119.830 ;
        RECT 0.805 118.385 7.195 118.675 ;
        RECT -2.215 116.470 -1.835 116.850 ;
        RECT 6.785 115.745 9.965 116.065 ;
      LAYER Metal2 ;
        RECT -2.885 119.490 -2.505 119.870 ;
        RECT -2.170 116.415 -1.870 123.455 ;
        RECT 0.855 118.285 1.175 123.445 ;
        RECT 6.865 115.685 7.145 118.720 ;
        RECT 9.615 115.640 9.915 122.795 ;
      LAYER Metal3 ;
        RECT -5.295 119.555 -2.500 119.850 ;
    END
  END b1_not
  PIN b1
    ANTENNADIFFAREA 2.559875 ;
    PORT
      LAYER Metal1 ;
        RECT 4.255 122.865 4.635 123.245 ;
        RECT 2.655 122.350 3.855 122.640 ;
        RECT -2.875 120.180 3.850 120.480 ;
        RECT 3.445 116.575 4.635 116.860 ;
        RECT 2.665 115.910 3.045 116.290 ;
      LAYER Metal2 ;
        RECT -2.850 120.160 -2.470 120.540 ;
        RECT 2.705 115.900 3.005 122.710 ;
        RECT 3.495 116.495 3.805 122.685 ;
        RECT 4.290 116.425 4.590 123.255 ;
      LAYER Metal3 ;
        RECT -5.330 120.185 -2.455 120.480 ;
    END
  END b1
  PIN a1_not_f
    ANTENNAGATEAREA 5.550000 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 29.575 125.100 31.030 125.480 ;
        RECT 29.735 122.800 31.030 123.180 ;
        RECT 43.220 122.800 44.530 123.180 ;
        RECT 28.065 121.475 44.075 121.850 ;
        RECT -2.895 120.895 10.665 121.195 ;
        RECT 12.570 120.895 30.990 121.195 ;
        RECT -0.430 117.220 2.490 117.520 ;
        RECT 6.035 117.205 9.405 117.505 ;
        RECT 15.030 117.220 17.950 117.520 ;
        RECT 21.495 117.205 24.865 117.505 ;
        RECT 29.745 117.300 31.050 117.680 ;
        RECT 43.085 117.300 44.550 117.680 ;
        RECT 29.560 115.300 31.050 115.680 ;
      LAYER Metal2 ;
        RECT -2.895 120.845 -2.515 121.225 ;
        RECT -0.395 117.170 -0.095 121.230 ;
        RECT 6.095 117.155 6.375 121.245 ;
        RECT 10.285 120.845 10.665 121.225 ;
        RECT 12.555 120.845 12.935 121.250 ;
        RECT 15.065 117.170 15.365 121.230 ;
        RECT 21.555 117.155 21.835 121.245 ;
        RECT 29.865 115.245 30.220 125.550 ;
        RECT 30.530 120.850 30.875 121.905 ;
        RECT 43.375 117.020 43.705 123.215 ;
      LAYER Metal3 ;
        RECT -5.335 120.900 -2.490 121.195 ;
        RECT 10.230 120.875 12.970 121.205 ;
    END
  END a1_not_f
  PIN a1_f
    ANTENNAGATEAREA 5.478500 ;
    ANTENNADIFFAREA 1.587600 ;
    PORT
      LAYER Metal1 ;
        RECT 53.270 125.200 54.550 125.580 ;
        RECT 39.770 122.800 40.955 123.180 ;
        RECT 53.270 122.800 54.285 123.180 ;
        RECT -2.890 121.640 10.675 121.955 ;
        RECT 12.565 121.640 26.390 121.940 ;
        RECT 28.065 120.120 54.295 120.510 ;
        RECT -1.660 118.985 2.470 119.285 ;
        RECT 4.845 118.935 9.345 119.245 ;
        RECT 13.800 118.985 17.930 119.285 ;
        RECT 20.305 118.935 24.805 119.245 ;
        RECT 39.750 117.300 41.110 117.680 ;
        RECT 53.250 117.300 54.430 117.680 ;
        RECT 53.250 115.300 54.325 115.680 ;
      LAYER Metal2 ;
        RECT -2.885 121.595 -2.505 121.975 ;
        RECT 10.280 121.595 10.660 121.975 ;
        RECT 12.550 121.595 12.930 122.000 ;
        RECT 26.015 121.595 26.375 123.425 ;
        RECT 28.195 120.075 28.610 123.425 ;
        RECT 40.390 123.165 40.700 123.195 ;
        RECT 40.390 117.065 40.705 123.165 ;
        RECT 53.890 115.070 54.220 125.765 ;
      LAYER Metal3 ;
        RECT 25.960 123.040 28.665 123.380 ;
        RECT -5.295 121.635 -2.470 121.940 ;
        RECT 10.225 121.625 12.970 121.955 ;
    END
  END a1_f
  OBS
      LAYER Nwell ;
        RECT -4.790 139.645 54.765 147.870 ;
      LAYER Pwell ;
        RECT -4.790 131.945 26.130 139.645 ;
        RECT 28.110 131.945 54.765 139.645 ;
      LAYER Nwell ;
        RECT 66.700 139.590 124.275 147.815 ;
      LAYER Pwell ;
        RECT 66.700 131.890 124.275 139.590 ;
      LAYER Nwell ;
        RECT -4.835 119.955 54.720 128.180 ;
      LAYER Pwell ;
        RECT -4.835 112.255 26.085 119.955 ;
        RECT 28.065 112.255 54.720 119.955 ;
      LAYER Nwell ;
        RECT 66.500 119.865 124.075 128.090 ;
      LAYER Pwell ;
        RECT 66.500 112.165 124.075 119.865 ;
      LAYER Nwell ;
        RECT -4.645 100.245 54.910 108.470 ;
      LAYER Pwell ;
        RECT -4.645 92.545 26.275 100.245 ;
        RECT 28.255 92.545 54.910 100.245 ;
      LAYER Nwell ;
        RECT 66.655 100.220 124.230 108.445 ;
      LAYER Pwell ;
        RECT 66.655 92.520 124.230 100.220 ;
      LAYER Nwell ;
        RECT -4.840 80.405 54.715 88.630 ;
      LAYER Pwell ;
        RECT -4.840 72.705 26.080 80.405 ;
        RECT 28.060 72.705 54.715 80.405 ;
      LAYER Nwell ;
        RECT 66.655 80.425 124.230 88.650 ;
      LAYER Pwell ;
        RECT 66.655 72.725 124.230 80.425 ;
      LAYER Nwell ;
        RECT -4.970 60.695 54.585 68.920 ;
      LAYER Pwell ;
        RECT -4.970 52.995 25.950 60.695 ;
        RECT 27.930 52.995 54.585 60.695 ;
      LAYER Nwell ;
        RECT 66.575 60.670 124.150 68.895 ;
      LAYER Pwell ;
        RECT 66.575 52.970 124.150 60.670 ;
      LAYER Nwell ;
        RECT -4.840 40.935 54.715 49.160 ;
      LAYER Pwell ;
        RECT -4.840 33.235 26.080 40.935 ;
        RECT 28.060 33.235 54.715 40.935 ;
      LAYER Nwell ;
        RECT 66.680 40.955 124.255 49.180 ;
      LAYER Pwell ;
        RECT 66.680 33.255 124.255 40.955 ;
      LAYER Nwell ;
        RECT -4.890 21.125 54.665 29.350 ;
      LAYER Pwell ;
        RECT -4.890 13.425 26.030 21.125 ;
        RECT 28.010 13.425 54.665 21.125 ;
      LAYER Nwell ;
        RECT 66.680 20.985 124.255 29.210 ;
      LAYER Pwell ;
        RECT 66.680 13.285 124.255 20.985 ;
      LAYER Nwell ;
        RECT -4.920 1.330 54.635 9.555 ;
      LAYER Pwell ;
        RECT -4.920 -6.370 26.000 1.330 ;
        RECT 27.980 -6.370 54.635 1.330 ;
      LAYER Nwell ;
        RECT 66.680 1.320 124.255 9.545 ;
      LAYER Pwell ;
        RECT 66.680 -6.380 124.255 1.320 ;
      LAYER Nwell ;
        RECT -4.770 -18.465 54.785 -10.240 ;
      LAYER Pwell ;
        RECT -4.770 -26.165 26.150 -18.465 ;
        RECT 28.130 -26.165 54.785 -18.465 ;
      LAYER Nwell ;
        RECT 66.720 -18.520 124.295 -10.295 ;
      LAYER Pwell ;
        RECT 66.720 -26.220 124.295 -18.520 ;
      LAYER Nwell ;
        RECT -4.815 -38.155 54.740 -29.930 ;
      LAYER Pwell ;
        RECT -4.815 -45.855 26.105 -38.155 ;
        RECT 28.085 -45.855 54.740 -38.155 ;
      LAYER Nwell ;
        RECT 66.520 -38.245 124.095 -30.020 ;
      LAYER Pwell ;
        RECT 66.520 -45.945 124.095 -38.245 ;
      LAYER Nwell ;
        RECT -4.625 -57.865 54.930 -49.640 ;
      LAYER Pwell ;
        RECT -4.625 -65.565 26.295 -57.865 ;
        RECT 28.275 -65.565 54.930 -57.865 ;
      LAYER Nwell ;
        RECT 66.675 -57.890 124.250 -49.665 ;
      LAYER Pwell ;
        RECT 66.675 -65.590 124.250 -57.890 ;
      LAYER Nwell ;
        RECT -4.820 -77.705 54.735 -69.480 ;
      LAYER Pwell ;
        RECT -4.820 -85.405 26.100 -77.705 ;
        RECT 28.080 -85.405 54.735 -77.705 ;
      LAYER Nwell ;
        RECT 66.675 -77.685 124.250 -69.460 ;
      LAYER Pwell ;
        RECT 66.675 -85.385 124.250 -77.685 ;
      LAYER Nwell ;
        RECT -4.950 -97.415 54.605 -89.190 ;
      LAYER Pwell ;
        RECT -4.950 -105.115 25.970 -97.415 ;
        RECT 27.950 -105.115 54.605 -97.415 ;
      LAYER Nwell ;
        RECT 66.595 -97.440 124.170 -89.215 ;
      LAYER Pwell ;
        RECT 66.595 -105.140 124.170 -97.440 ;
      LAYER Nwell ;
        RECT -4.820 -117.175 54.735 -108.950 ;
      LAYER Pwell ;
        RECT -4.820 -124.875 26.100 -117.175 ;
        RECT 28.080 -124.875 54.735 -117.175 ;
      LAYER Nwell ;
        RECT 66.700 -117.155 124.275 -108.930 ;
      LAYER Pwell ;
        RECT 66.700 -124.855 124.275 -117.155 ;
      LAYER Nwell ;
        RECT -4.870 -136.985 54.685 -128.760 ;
      LAYER Pwell ;
        RECT -4.870 -144.685 26.050 -136.985 ;
        RECT 28.030 -144.685 54.685 -136.985 ;
      LAYER Nwell ;
        RECT 66.700 -137.125 124.275 -128.900 ;
      LAYER Pwell ;
        RECT 66.700 -144.825 124.275 -137.125 ;
      LAYER Nwell ;
        RECT -4.900 -156.780 54.655 -148.555 ;
      LAYER Pwell ;
        RECT -4.900 -164.480 26.020 -156.780 ;
        RECT 28.000 -164.480 54.655 -156.780 ;
      LAYER Nwell ;
        RECT 66.700 -156.790 124.275 -148.565 ;
      LAYER Pwell ;
        RECT 66.700 -164.490 124.275 -156.790 ;
      LAYER Metal1 ;
        RECT -4.360 147.815 68.030 147.870 ;
        RECT -4.360 146.970 124.275 147.815 ;
        RECT -3.990 139.810 -3.610 146.970 ;
        RECT 1.585 142.515 1.965 142.895 ;
        RECT 8.485 142.505 8.865 142.885 ;
        RECT -1.090 142.090 0.650 142.380 ;
        RECT 5.410 142.010 8.020 142.435 ;
        RECT 7.595 139.570 10.700 139.845 ;
        RECT 11.470 139.810 11.850 146.970 ;
        RECT 67.920 146.915 124.275 146.970 ;
        RECT 28.110 145.930 65.660 145.985 ;
        RECT 28.110 145.700 93.680 145.930 ;
        RECT 64.905 145.645 93.680 145.700 ;
        RECT 95.350 145.625 102.055 145.925 ;
        RECT 31.815 144.790 33.015 145.170 ;
        RECT 34.770 144.575 37.045 145.085 ;
        RECT 39.670 144.575 41.970 145.085 ;
        RECT 44.265 144.575 46.545 145.085 ;
        RECT 51.340 144.890 52.575 145.270 ;
        RECT 68.210 144.735 69.665 145.115 ;
        RECT 52.755 144.535 53.135 144.570 ;
        RECT 31.255 144.430 31.635 144.470 ;
        RECT 31.185 144.125 34.020 144.430 ;
        RECT 50.000 144.225 53.135 144.535 ;
        RECT 73.360 144.520 75.635 145.030 ;
        RECT 78.260 144.520 80.560 145.030 ;
        RECT 82.855 144.520 85.135 145.030 ;
        RECT 91.905 144.835 93.185 145.215 ;
        RECT 91.345 144.480 91.725 144.515 ;
        RECT 69.845 144.375 70.225 144.415 ;
        RECT 52.755 144.190 53.135 144.225 ;
        RECT 31.255 144.090 31.635 144.125 ;
        RECT 69.775 144.070 72.610 144.375 ;
        RECT 88.590 144.170 91.725 144.480 ;
        RECT 91.345 144.135 91.725 144.170 ;
        RECT 69.845 144.035 70.225 144.070 ;
        RECT 13.300 142.715 16.705 143.155 ;
        RECT 17.045 142.515 17.425 142.895 ;
        RECT 19.760 142.555 20.140 142.935 ;
        RECT 23.945 142.505 24.325 142.885 ;
        RECT 31.815 142.490 35.075 142.870 ;
        RECT 35.815 142.490 39.075 142.870 ;
        RECT 45.315 142.490 48.575 142.870 ;
        RECT 49.315 142.490 52.575 142.870 ;
        RECT 14.370 142.090 16.110 142.380 ;
        RECT 18.160 142.040 19.360 142.330 ;
        RECT 20.870 142.010 23.465 142.385 ;
        RECT 25.080 142.105 25.460 142.485 ;
        RECT 68.370 142.435 69.665 142.815 ;
        RECT 74.405 142.435 77.665 142.815 ;
        RECT 78.405 142.435 79.590 142.815 ;
        RECT 81.855 142.435 83.165 142.815 ;
        RECT 83.905 142.435 87.165 142.815 ;
        RECT 91.905 142.435 92.920 142.815 ;
        RECT 95.985 142.680 99.400 143.100 ;
        RECT 99.730 142.460 100.110 142.840 ;
        RECT 102.445 142.500 102.825 142.880 ;
        RECT 106.630 142.450 107.010 142.830 ;
        RECT 31.255 141.790 31.635 142.170 ;
        RECT 35.255 141.790 35.635 142.170 ;
        RECT 39.255 142.125 39.635 142.170 ;
        RECT 44.755 142.125 45.135 142.170 ;
        RECT 39.205 141.810 45.140 142.125 ;
        RECT 39.255 141.790 39.635 141.810 ;
        RECT 44.755 141.790 45.135 141.810 ;
        RECT 48.755 141.790 49.135 142.170 ;
        RECT 52.755 141.790 53.135 142.170 ;
        RECT 69.845 141.735 70.225 142.115 ;
        RECT 73.845 141.735 74.225 142.115 ;
        RECT 77.845 142.070 78.225 142.115 ;
        RECT 83.345 142.070 83.725 142.115 ;
        RECT 77.795 141.755 83.730 142.070 ;
        RECT 77.845 141.735 78.225 141.755 ;
        RECT 83.345 141.735 83.725 141.755 ;
        RECT 87.345 141.735 87.725 142.115 ;
        RECT 91.345 141.735 91.725 142.115 ;
        RECT 97.055 142.035 98.795 142.325 ;
        RECT 100.845 141.985 102.045 142.275 ;
        RECT 103.555 141.945 106.185 142.400 ;
        RECT 107.765 142.050 108.145 142.430 ;
        RECT 61.935 141.110 82.710 141.485 ;
        RECT 32.480 140.575 59.790 140.915 ;
        RECT 12.095 139.870 19.355 140.170 ;
        RECT 12.650 139.335 16.735 139.605 ;
        RECT 23.055 139.570 26.805 139.845 ;
        RECT 60.965 139.755 92.930 140.145 ;
        RECT 105.740 139.515 108.870 139.790 ;
        RECT 109.615 139.755 109.995 146.915 ;
        RECT 110.855 144.455 117.595 144.755 ;
        RECT 111.445 142.660 114.900 143.100 ;
        RECT 117.905 142.500 118.285 142.880 ;
        RECT 116.305 141.985 117.505 142.275 ;
        RECT 123.225 142.050 123.605 142.430 ;
        RECT 110.260 141.275 126.180 141.575 ;
        RECT 110.795 140.530 127.740 140.830 ;
        RECT 28.110 139.445 46.780 139.455 ;
        RECT 28.110 139.400 58.130 139.445 ;
        RECT 28.110 139.390 85.370 139.400 ;
        RECT 28.110 139.135 94.375 139.390 ;
        RECT 57.810 139.080 94.375 139.135 ;
        RECT -3.990 132.845 -3.610 138.675 ;
        RECT 0.265 137.495 10.920 137.830 ;
        RECT 0.235 136.175 2.015 136.465 ;
        RECT 7.610 136.145 8.920 136.465 ;
        RECT -1.035 135.560 -0.655 135.940 ;
        RECT 5.420 135.590 5.800 135.970 ;
        RECT -3.240 132.845 0.855 132.850 ;
        RECT 11.470 132.845 11.850 138.675 ;
        RECT 111.990 138.620 116.120 138.920 ;
        RECT 27.580 138.410 63.490 138.465 ;
        RECT 16.310 138.075 22.700 138.365 ;
        RECT 27.580 138.195 94.775 138.410 ;
        RECT 63.030 138.140 94.775 138.195 ;
        RECT 98.995 138.020 105.385 138.310 ;
        RECT 15.725 137.495 26.230 137.830 ;
        RECT 51.200 137.630 61.750 137.965 ;
        RECT 98.410 137.440 108.890 137.775 ;
        RECT 31.795 136.990 35.095 137.370 ;
        RECT 35.795 136.990 39.095 137.370 ;
        RECT 45.295 136.990 48.595 137.370 ;
        RECT 49.295 136.990 52.595 137.370 ;
        RECT 68.380 136.935 69.685 137.315 ;
        RECT 74.385 136.935 77.685 137.315 ;
        RECT 78.385 136.935 79.745 137.315 ;
        RECT 81.720 136.935 83.185 137.315 ;
        RECT 83.885 136.935 87.185 137.315 ;
        RECT 91.885 136.935 93.065 137.315 ;
        RECT 31.255 136.645 31.635 136.680 ;
        RECT 13.290 136.160 13.670 136.540 ;
        RECT 15.695 136.175 17.475 136.465 ;
        RECT 18.950 136.265 20.140 136.550 ;
        RECT 23.070 136.145 24.380 136.465 ;
        RECT 30.990 136.335 34.000 136.645 ;
        RECT 31.255 136.300 31.635 136.335 ;
        RECT 35.255 136.300 36.345 136.680 ;
        RECT 39.255 136.675 39.635 136.680 ;
        RECT 36.775 136.310 39.640 136.675 ;
        RECT 44.755 136.655 45.135 136.680 ;
        RECT 44.740 136.335 46.885 136.655 ;
        RECT 39.255 136.300 39.635 136.310 ;
        RECT 44.755 136.300 45.135 136.335 ;
        RECT 47.800 136.300 49.135 136.680 ;
        RECT 52.755 136.660 53.135 136.680 ;
        RECT 50.290 136.340 53.200 136.660 ;
        RECT 69.845 136.590 70.225 136.625 ;
        RECT 52.755 136.300 53.135 136.340 ;
        RECT 69.580 136.280 72.590 136.590 ;
        RECT 69.845 136.245 70.225 136.280 ;
        RECT 73.845 136.245 74.935 136.625 ;
        RECT 77.845 136.620 78.225 136.625 ;
        RECT 75.365 136.255 78.230 136.620 ;
        RECT 83.345 136.600 83.725 136.625 ;
        RECT 83.330 136.280 85.475 136.600 ;
        RECT 77.845 136.245 78.225 136.255 ;
        RECT 83.345 136.245 83.725 136.280 ;
        RECT 86.390 136.245 87.725 136.625 ;
        RECT 91.345 136.605 91.725 136.625 ;
        RECT 88.880 136.285 91.790 136.605 ;
        RECT 91.345 136.245 91.725 136.285 ;
        RECT 95.975 136.105 96.355 136.485 ;
        RECT 98.380 136.120 100.160 136.410 ;
        RECT 101.635 136.210 102.825 136.495 ;
        RECT 105.755 136.090 107.065 136.410 ;
        RECT 14.425 135.560 14.805 135.940 ;
        RECT 18.170 135.600 18.550 135.980 ;
        RECT 20.880 135.590 21.260 135.970 ;
        RECT 22.290 135.435 25.470 135.755 ;
        RECT 97.110 135.505 97.490 135.885 ;
        RECT 100.855 135.545 101.235 135.925 ;
        RECT 103.565 135.535 103.945 135.915 ;
        RECT 104.975 135.380 108.155 135.700 ;
        RECT 31.795 134.990 33.080 135.370 ;
        RECT 51.110 134.990 52.595 135.370 ;
        RECT 68.195 134.935 69.685 135.315 ;
        RECT 91.885 134.935 92.960 135.315 ;
        RECT 31.255 134.300 32.345 134.680 ;
        RECT 33.300 134.310 34.820 134.670 ;
        RECT 35.740 134.305 48.590 134.640 ;
        RECT 52.755 134.635 53.135 134.680 ;
        RECT 52.020 134.335 53.330 134.635 ;
        RECT 52.755 134.300 53.135 134.335 ;
        RECT 69.845 134.245 70.935 134.625 ;
        RECT 71.890 134.255 73.410 134.615 ;
        RECT 74.330 134.250 87.180 134.585 ;
        RECT 91.345 134.580 91.725 134.625 ;
        RECT 90.610 134.280 91.920 134.580 ;
        RECT 91.345 134.245 91.725 134.280 ;
        RECT 28.110 133.750 61.190 133.790 ;
        RECT 28.110 133.440 93.355 133.750 ;
        RECT 60.405 133.385 93.355 133.440 ;
        RECT 95.150 133.375 99.410 133.730 ;
        RECT 12.220 132.845 16.315 132.850 ;
        RECT -4.360 132.840 0.855 132.845 ;
        RECT 11.100 132.840 16.315 132.845 ;
        RECT 26.560 132.840 66.810 132.845 ;
        RECT -4.360 132.790 66.810 132.840 ;
        RECT 93.355 132.790 99.000 132.795 ;
        RECT 109.615 132.790 109.995 138.620 ;
        RECT 118.495 138.570 122.995 138.880 ;
        RECT 114.455 138.020 120.845 138.310 ;
        RECT 113.220 136.855 116.140 137.155 ;
        RECT 119.685 136.840 123.055 137.140 ;
        RECT 111.435 136.105 111.815 136.485 ;
        RECT 117.095 136.210 118.285 136.495 ;
        RECT 116.315 135.545 116.695 135.925 ;
        RECT 120.435 135.380 123.615 135.700 ;
        RECT 110.715 134.295 114.865 134.565 ;
        RECT 110.365 132.790 114.460 132.795 ;
        RECT -4.360 132.785 99.000 132.790 ;
        RECT 109.245 132.785 114.460 132.790 ;
        RECT -4.360 131.945 124.275 132.785 ;
        RECT 66.700 131.890 124.275 131.945 ;
        RECT -4.405 128.090 67.985 128.180 ;
        RECT -4.405 127.280 124.075 128.090 ;
        RECT -4.035 120.120 -3.655 127.280 ;
        RECT 1.540 122.825 1.920 123.205 ;
        RECT 8.440 122.815 8.820 123.195 ;
        RECT -1.135 122.400 0.605 122.690 ;
        RECT 5.365 122.320 7.975 122.745 ;
        RECT 7.550 119.880 10.655 120.155 ;
        RECT 11.425 120.120 11.805 127.280 ;
        RECT 67.720 127.190 124.075 127.280 ;
        RECT 28.065 126.205 65.615 126.295 ;
        RECT 28.065 126.010 93.480 126.205 ;
        RECT 64.705 125.920 93.480 126.010 ;
        RECT 95.150 125.900 101.855 126.200 ;
        RECT 31.770 125.100 32.970 125.480 ;
        RECT 34.725 124.885 37.000 125.395 ;
        RECT 39.625 124.885 41.925 125.395 ;
        RECT 44.220 124.885 46.500 125.395 ;
        RECT 51.295 125.200 52.530 125.580 ;
        RECT 68.010 125.010 69.465 125.390 ;
        RECT 52.710 124.845 53.090 124.880 ;
        RECT 31.210 124.740 31.590 124.780 ;
        RECT 31.140 124.435 33.975 124.740 ;
        RECT 49.955 124.535 53.090 124.845 ;
        RECT 73.160 124.795 75.435 125.305 ;
        RECT 78.060 124.795 80.360 125.305 ;
        RECT 82.655 124.795 84.935 125.305 ;
        RECT 91.705 125.110 92.985 125.490 ;
        RECT 91.145 124.755 91.525 124.790 ;
        RECT 69.645 124.650 70.025 124.690 ;
        RECT 52.710 124.500 53.090 124.535 ;
        RECT 31.210 124.400 31.590 124.435 ;
        RECT 69.575 124.345 72.410 124.650 ;
        RECT 88.390 124.445 91.525 124.755 ;
        RECT 91.145 124.410 91.525 124.445 ;
        RECT 69.645 124.310 70.025 124.345 ;
        RECT 13.255 123.025 16.660 123.465 ;
        RECT 17.000 122.825 17.380 123.205 ;
        RECT 19.715 122.865 20.095 123.245 ;
        RECT 23.900 122.815 24.280 123.195 ;
        RECT 31.770 122.800 35.030 123.180 ;
        RECT 35.770 122.800 39.030 123.180 ;
        RECT 45.270 122.800 48.530 123.180 ;
        RECT 49.270 122.800 52.530 123.180 ;
        RECT 14.325 122.400 16.065 122.690 ;
        RECT 18.115 122.350 19.315 122.640 ;
        RECT 20.825 122.320 23.420 122.695 ;
        RECT 25.035 122.415 25.415 122.795 ;
        RECT 68.170 122.710 69.465 123.090 ;
        RECT 74.205 122.710 77.465 123.090 ;
        RECT 78.205 122.710 79.390 123.090 ;
        RECT 81.655 122.710 82.965 123.090 ;
        RECT 83.705 122.710 86.965 123.090 ;
        RECT 91.705 122.710 92.720 123.090 ;
        RECT 95.785 122.955 99.200 123.375 ;
        RECT 99.530 122.735 99.910 123.115 ;
        RECT 102.245 122.775 102.625 123.155 ;
        RECT 106.430 122.725 106.810 123.105 ;
        RECT 31.210 122.100 31.590 122.480 ;
        RECT 35.210 122.100 35.590 122.480 ;
        RECT 39.210 122.435 39.590 122.480 ;
        RECT 44.710 122.435 45.090 122.480 ;
        RECT 39.160 122.120 45.095 122.435 ;
        RECT 39.210 122.100 39.590 122.120 ;
        RECT 44.710 122.100 45.090 122.120 ;
        RECT 48.710 122.100 49.090 122.480 ;
        RECT 52.710 122.100 53.090 122.480 ;
        RECT 69.645 122.010 70.025 122.390 ;
        RECT 73.645 122.010 74.025 122.390 ;
        RECT 77.645 122.345 78.025 122.390 ;
        RECT 83.145 122.345 83.525 122.390 ;
        RECT 77.595 122.030 83.530 122.345 ;
        RECT 77.645 122.010 78.025 122.030 ;
        RECT 83.145 122.010 83.525 122.030 ;
        RECT 87.145 122.010 87.525 122.390 ;
        RECT 91.145 122.010 91.525 122.390 ;
        RECT 96.855 122.310 98.595 122.600 ;
        RECT 100.645 122.260 101.845 122.550 ;
        RECT 103.355 122.220 105.985 122.675 ;
        RECT 107.565 122.325 107.945 122.705 ;
        RECT 61.735 121.385 82.510 121.760 ;
        RECT 32.435 120.885 59.745 121.225 ;
        RECT 12.050 120.180 19.310 120.480 ;
        RECT 12.605 119.645 16.690 119.915 ;
        RECT 23.010 119.880 26.760 120.155 ;
        RECT 60.765 120.030 92.730 120.420 ;
        RECT 105.540 119.790 108.670 120.065 ;
        RECT 109.415 120.030 109.795 127.190 ;
        RECT 110.655 124.730 117.395 125.030 ;
        RECT 111.245 122.935 114.700 123.375 ;
        RECT 117.705 122.775 118.085 123.155 ;
        RECT 116.105 122.260 117.305 122.550 ;
        RECT 123.025 122.325 123.405 122.705 ;
        RECT 110.060 121.550 125.980 121.850 ;
        RECT 110.595 120.805 127.540 121.105 ;
        RECT 28.065 119.755 46.735 119.765 ;
        RECT 28.065 119.675 58.085 119.755 ;
        RECT 28.065 119.665 85.170 119.675 ;
        RECT 28.065 119.445 94.175 119.665 ;
        RECT 57.610 119.355 94.175 119.445 ;
        RECT -4.035 113.155 -3.655 118.985 ;
        RECT 0.220 117.805 10.875 118.140 ;
        RECT 0.190 116.485 1.970 116.775 ;
        RECT 7.565 116.455 8.875 116.775 ;
        RECT -1.080 115.870 -0.700 116.250 ;
        RECT 5.375 115.900 5.755 116.280 ;
        RECT -3.285 113.155 0.810 113.160 ;
        RECT 11.425 113.155 11.805 118.985 ;
        RECT 111.790 118.895 115.920 119.195 ;
        RECT 27.535 118.685 63.445 118.775 ;
        RECT 16.265 118.385 22.655 118.675 ;
        RECT 27.535 118.505 94.575 118.685 ;
        RECT 62.830 118.415 94.575 118.505 ;
        RECT 98.795 118.295 105.185 118.585 ;
        RECT 15.680 117.805 26.185 118.140 ;
        RECT 51.155 117.940 61.705 118.275 ;
        RECT 98.210 117.715 108.690 118.050 ;
        RECT 31.750 117.300 35.050 117.680 ;
        RECT 35.750 117.300 39.050 117.680 ;
        RECT 45.250 117.300 48.550 117.680 ;
        RECT 49.250 117.300 52.550 117.680 ;
        RECT 68.180 117.210 69.485 117.590 ;
        RECT 74.185 117.210 77.485 117.590 ;
        RECT 78.185 117.210 79.545 117.590 ;
        RECT 81.520 117.210 82.985 117.590 ;
        RECT 83.685 117.210 86.985 117.590 ;
        RECT 91.685 117.210 92.865 117.590 ;
        RECT 31.210 116.955 31.590 116.990 ;
        RECT 13.245 116.470 13.625 116.850 ;
        RECT 15.650 116.485 17.430 116.775 ;
        RECT 18.905 116.575 20.095 116.860 ;
        RECT 23.025 116.455 24.335 116.775 ;
        RECT 30.945 116.645 33.955 116.955 ;
        RECT 31.210 116.610 31.590 116.645 ;
        RECT 35.210 116.610 36.300 116.990 ;
        RECT 39.210 116.985 39.590 116.990 ;
        RECT 36.730 116.620 39.595 116.985 ;
        RECT 44.710 116.965 45.090 116.990 ;
        RECT 44.695 116.645 46.840 116.965 ;
        RECT 39.210 116.610 39.590 116.620 ;
        RECT 44.710 116.610 45.090 116.645 ;
        RECT 47.755 116.610 49.090 116.990 ;
        RECT 52.710 116.970 53.090 116.990 ;
        RECT 50.245 116.650 53.155 116.970 ;
        RECT 69.645 116.865 70.025 116.900 ;
        RECT 52.710 116.610 53.090 116.650 ;
        RECT 69.380 116.555 72.390 116.865 ;
        RECT 69.645 116.520 70.025 116.555 ;
        RECT 73.645 116.520 74.735 116.900 ;
        RECT 77.645 116.895 78.025 116.900 ;
        RECT 75.165 116.530 78.030 116.895 ;
        RECT 83.145 116.875 83.525 116.900 ;
        RECT 83.130 116.555 85.275 116.875 ;
        RECT 77.645 116.520 78.025 116.530 ;
        RECT 83.145 116.520 83.525 116.555 ;
        RECT 86.190 116.520 87.525 116.900 ;
        RECT 91.145 116.880 91.525 116.900 ;
        RECT 88.680 116.560 91.590 116.880 ;
        RECT 91.145 116.520 91.525 116.560 ;
        RECT 95.775 116.380 96.155 116.760 ;
        RECT 98.180 116.395 99.960 116.685 ;
        RECT 101.435 116.485 102.625 116.770 ;
        RECT 105.555 116.365 106.865 116.685 ;
        RECT 14.380 115.870 14.760 116.250 ;
        RECT 18.125 115.910 18.505 116.290 ;
        RECT 20.835 115.900 21.215 116.280 ;
        RECT 22.245 115.745 25.425 116.065 ;
        RECT 96.910 115.780 97.290 116.160 ;
        RECT 100.655 115.820 101.035 116.200 ;
        RECT 103.365 115.810 103.745 116.190 ;
        RECT 31.750 115.300 33.035 115.680 ;
        RECT 51.065 115.300 52.550 115.680 ;
        RECT 104.775 115.655 107.955 115.975 ;
        RECT 67.995 115.210 69.485 115.590 ;
        RECT 91.685 115.210 92.760 115.590 ;
        RECT 31.210 114.610 32.300 114.990 ;
        RECT 33.255 114.620 34.775 114.980 ;
        RECT 35.695 114.615 48.545 114.950 ;
        RECT 52.710 114.945 53.090 114.990 ;
        RECT 51.975 114.645 53.285 114.945 ;
        RECT 52.710 114.610 53.090 114.645 ;
        RECT 69.645 114.520 70.735 114.900 ;
        RECT 71.690 114.530 73.210 114.890 ;
        RECT 74.130 114.525 86.980 114.860 ;
        RECT 91.145 114.855 91.525 114.900 ;
        RECT 90.410 114.555 91.720 114.855 ;
        RECT 91.145 114.520 91.525 114.555 ;
        RECT 28.065 114.025 61.145 114.100 ;
        RECT 28.065 113.750 93.155 114.025 ;
        RECT 60.205 113.660 93.155 113.750 ;
        RECT 94.950 113.650 99.210 114.005 ;
        RECT 12.175 113.155 16.270 113.160 ;
        RECT -4.405 113.150 0.810 113.155 ;
        RECT 11.055 113.150 16.270 113.155 ;
        RECT 26.515 113.150 66.765 113.155 ;
        RECT -4.405 113.065 66.765 113.150 ;
        RECT 93.155 113.065 98.800 113.070 ;
        RECT 109.415 113.065 109.795 118.895 ;
        RECT 118.295 118.845 122.795 119.155 ;
        RECT 114.255 118.295 120.645 118.585 ;
        RECT 113.020 117.130 115.940 117.430 ;
        RECT 119.485 117.115 122.855 117.415 ;
        RECT 111.235 116.380 111.615 116.760 ;
        RECT 116.895 116.485 118.085 116.770 ;
        RECT 116.115 115.820 116.495 116.200 ;
        RECT 120.235 115.655 123.415 115.975 ;
        RECT 110.515 114.570 114.665 114.840 ;
        RECT 110.165 113.065 114.260 113.070 ;
        RECT -4.405 113.060 98.800 113.065 ;
        RECT 109.045 113.060 114.260 113.065 ;
        RECT -4.405 112.255 124.075 113.060 ;
        RECT 66.500 112.165 124.075 112.255 ;
        RECT -4.215 108.445 68.175 108.470 ;
        RECT -4.215 107.570 124.230 108.445 ;
        RECT -3.845 100.410 -3.465 107.570 ;
        RECT 1.730 103.115 2.110 103.495 ;
        RECT 8.630 103.105 9.010 103.485 ;
        RECT -0.945 102.690 0.795 102.980 ;
        RECT 5.555 102.610 8.165 103.035 ;
        RECT 7.740 100.170 10.845 100.445 ;
        RECT 11.615 100.410 11.995 107.570 ;
        RECT 67.875 107.545 124.230 107.570 ;
        RECT 28.255 106.560 65.805 106.585 ;
        RECT 28.255 106.300 93.635 106.560 ;
        RECT 64.860 106.275 93.635 106.300 ;
        RECT 95.305 106.255 102.010 106.555 ;
        RECT 31.960 105.390 33.160 105.770 ;
        RECT 34.915 105.175 37.190 105.685 ;
        RECT 39.815 105.175 42.115 105.685 ;
        RECT 44.410 105.175 46.690 105.685 ;
        RECT 51.485 105.490 52.720 105.870 ;
        RECT 68.165 105.365 69.620 105.745 ;
        RECT 52.900 105.135 53.280 105.170 ;
        RECT 73.315 105.150 75.590 105.660 ;
        RECT 78.215 105.150 80.515 105.660 ;
        RECT 82.810 105.150 85.090 105.660 ;
        RECT 91.860 105.465 93.140 105.845 ;
        RECT 31.400 105.030 31.780 105.070 ;
        RECT 31.330 104.725 34.165 105.030 ;
        RECT 50.145 104.825 53.280 105.135 ;
        RECT 91.300 105.110 91.680 105.145 ;
        RECT 69.800 105.005 70.180 105.045 ;
        RECT 52.900 104.790 53.280 104.825 ;
        RECT 31.400 104.690 31.780 104.725 ;
        RECT 69.730 104.700 72.565 105.005 ;
        RECT 88.545 104.800 91.680 105.110 ;
        RECT 91.300 104.765 91.680 104.800 ;
        RECT 69.800 104.665 70.180 104.700 ;
        RECT 13.445 103.315 16.850 103.755 ;
        RECT 17.190 103.115 17.570 103.495 ;
        RECT 19.905 103.155 20.285 103.535 ;
        RECT 24.090 103.105 24.470 103.485 ;
        RECT 31.960 103.090 35.220 103.470 ;
        RECT 35.960 103.090 39.220 103.470 ;
        RECT 45.460 103.090 48.720 103.470 ;
        RECT 49.460 103.090 52.720 103.470 ;
        RECT 14.515 102.690 16.255 102.980 ;
        RECT 18.305 102.640 19.505 102.930 ;
        RECT 21.015 102.610 23.610 102.985 ;
        RECT 25.225 102.705 25.605 103.085 ;
        RECT 68.325 103.065 69.620 103.445 ;
        RECT 74.360 103.065 77.620 103.445 ;
        RECT 78.360 103.065 79.545 103.445 ;
        RECT 81.810 103.065 83.120 103.445 ;
        RECT 83.860 103.065 87.120 103.445 ;
        RECT 91.860 103.065 92.875 103.445 ;
        RECT 95.940 103.310 99.355 103.730 ;
        RECT 99.685 103.090 100.065 103.470 ;
        RECT 102.400 103.130 102.780 103.510 ;
        RECT 106.585 103.080 106.965 103.460 ;
        RECT 31.400 102.390 31.780 102.770 ;
        RECT 35.400 102.390 35.780 102.770 ;
        RECT 39.400 102.725 39.780 102.770 ;
        RECT 44.900 102.725 45.280 102.770 ;
        RECT 39.350 102.410 45.285 102.725 ;
        RECT 39.400 102.390 39.780 102.410 ;
        RECT 44.900 102.390 45.280 102.410 ;
        RECT 48.900 102.390 49.280 102.770 ;
        RECT 52.900 102.390 53.280 102.770 ;
        RECT 69.800 102.365 70.180 102.745 ;
        RECT 73.800 102.365 74.180 102.745 ;
        RECT 77.800 102.700 78.180 102.745 ;
        RECT 83.300 102.700 83.680 102.745 ;
        RECT 77.750 102.385 83.685 102.700 ;
        RECT 77.800 102.365 78.180 102.385 ;
        RECT 83.300 102.365 83.680 102.385 ;
        RECT 87.300 102.365 87.680 102.745 ;
        RECT 91.300 102.365 91.680 102.745 ;
        RECT 97.010 102.665 98.750 102.955 ;
        RECT 100.800 102.615 102.000 102.905 ;
        RECT 103.510 102.575 106.140 103.030 ;
        RECT 107.720 102.680 108.100 103.060 ;
        RECT 61.890 101.740 82.665 102.115 ;
        RECT 32.625 101.175 59.935 101.515 ;
        RECT 12.240 100.470 19.500 100.770 ;
        RECT 12.795 99.935 16.880 100.205 ;
        RECT 23.200 100.170 26.950 100.445 ;
        RECT 60.920 100.385 92.885 100.775 ;
        RECT 105.695 100.145 108.825 100.420 ;
        RECT 109.570 100.385 109.950 107.545 ;
        RECT 110.810 105.085 117.550 105.385 ;
        RECT 111.400 103.290 114.855 103.730 ;
        RECT 117.860 103.130 118.240 103.510 ;
        RECT 116.260 102.615 117.460 102.905 ;
        RECT 123.180 102.680 123.560 103.060 ;
        RECT 110.215 101.905 126.135 102.205 ;
        RECT 110.750 101.160 127.695 101.460 ;
        RECT 28.255 100.045 46.925 100.055 ;
        RECT 28.255 100.030 58.275 100.045 ;
        RECT 28.255 100.020 85.325 100.030 ;
        RECT 28.255 99.735 94.330 100.020 ;
        RECT 57.765 99.710 94.330 99.735 ;
        RECT -3.845 93.445 -3.465 99.275 ;
        RECT 0.410 98.095 11.065 98.430 ;
        RECT 0.380 96.775 2.160 97.065 ;
        RECT 7.755 96.745 9.065 97.065 ;
        RECT -0.890 96.160 -0.510 96.540 ;
        RECT 5.565 96.190 5.945 96.570 ;
        RECT -3.095 93.445 1.000 93.450 ;
        RECT 11.615 93.445 11.995 99.275 ;
        RECT 111.945 99.250 116.075 99.550 ;
        RECT 27.725 99.040 63.635 99.065 ;
        RECT 16.455 98.675 22.845 98.965 ;
        RECT 27.725 98.795 94.730 99.040 ;
        RECT 62.985 98.770 94.730 98.795 ;
        RECT 98.950 98.650 105.340 98.940 ;
        RECT 15.870 98.095 26.375 98.430 ;
        RECT 51.345 98.230 61.895 98.565 ;
        RECT 98.365 98.070 108.845 98.405 ;
        RECT 31.940 97.590 35.240 97.970 ;
        RECT 35.940 97.590 39.240 97.970 ;
        RECT 45.440 97.590 48.740 97.970 ;
        RECT 49.440 97.590 52.740 97.970 ;
        RECT 68.335 97.565 69.640 97.945 ;
        RECT 74.340 97.565 77.640 97.945 ;
        RECT 78.340 97.565 79.700 97.945 ;
        RECT 81.675 97.565 83.140 97.945 ;
        RECT 83.840 97.565 87.140 97.945 ;
        RECT 91.840 97.565 93.020 97.945 ;
        RECT 31.400 97.245 31.780 97.280 ;
        RECT 13.435 96.760 13.815 97.140 ;
        RECT 15.840 96.775 17.620 97.065 ;
        RECT 19.095 96.865 20.285 97.150 ;
        RECT 23.215 96.745 24.525 97.065 ;
        RECT 31.135 96.935 34.145 97.245 ;
        RECT 31.400 96.900 31.780 96.935 ;
        RECT 35.400 96.900 36.490 97.280 ;
        RECT 39.400 97.275 39.780 97.280 ;
        RECT 36.920 96.910 39.785 97.275 ;
        RECT 44.900 97.255 45.280 97.280 ;
        RECT 44.885 96.935 47.030 97.255 ;
        RECT 39.400 96.900 39.780 96.910 ;
        RECT 44.900 96.900 45.280 96.935 ;
        RECT 47.945 96.900 49.280 97.280 ;
        RECT 52.900 97.260 53.280 97.280 ;
        RECT 50.435 96.940 53.345 97.260 ;
        RECT 69.800 97.220 70.180 97.255 ;
        RECT 52.900 96.900 53.280 96.940 ;
        RECT 69.535 96.910 72.545 97.220 ;
        RECT 69.800 96.875 70.180 96.910 ;
        RECT 73.800 96.875 74.890 97.255 ;
        RECT 77.800 97.250 78.180 97.255 ;
        RECT 75.320 96.885 78.185 97.250 ;
        RECT 83.300 97.230 83.680 97.255 ;
        RECT 83.285 96.910 85.430 97.230 ;
        RECT 77.800 96.875 78.180 96.885 ;
        RECT 83.300 96.875 83.680 96.910 ;
        RECT 86.345 96.875 87.680 97.255 ;
        RECT 91.300 97.235 91.680 97.255 ;
        RECT 88.835 96.915 91.745 97.235 ;
        RECT 91.300 96.875 91.680 96.915 ;
        RECT 95.930 96.735 96.310 97.115 ;
        RECT 98.335 96.750 100.115 97.040 ;
        RECT 101.590 96.840 102.780 97.125 ;
        RECT 105.710 96.720 107.020 97.040 ;
        RECT 14.570 96.160 14.950 96.540 ;
        RECT 18.315 96.200 18.695 96.580 ;
        RECT 21.025 96.190 21.405 96.570 ;
        RECT 22.435 96.035 25.615 96.355 ;
        RECT 97.065 96.135 97.445 96.515 ;
        RECT 100.810 96.175 101.190 96.555 ;
        RECT 103.520 96.165 103.900 96.545 ;
        RECT 104.930 96.010 108.110 96.330 ;
        RECT 31.940 95.590 33.225 95.970 ;
        RECT 51.255 95.590 52.740 95.970 ;
        RECT 68.150 95.565 69.640 95.945 ;
        RECT 91.840 95.565 92.915 95.945 ;
        RECT 31.400 94.900 32.490 95.280 ;
        RECT 33.445 94.910 34.965 95.270 ;
        RECT 35.885 94.905 48.735 95.240 ;
        RECT 52.900 95.235 53.280 95.280 ;
        RECT 52.165 94.935 53.475 95.235 ;
        RECT 52.900 94.900 53.280 94.935 ;
        RECT 69.800 94.875 70.890 95.255 ;
        RECT 71.845 94.885 73.365 95.245 ;
        RECT 74.285 94.880 87.135 95.215 ;
        RECT 91.300 95.210 91.680 95.255 ;
        RECT 90.565 94.910 91.875 95.210 ;
        RECT 91.300 94.875 91.680 94.910 ;
        RECT 28.255 94.380 61.335 94.390 ;
        RECT 28.255 94.040 93.310 94.380 ;
        RECT 60.360 94.015 93.310 94.040 ;
        RECT 95.105 94.005 99.365 94.360 ;
        RECT 12.365 93.445 16.460 93.450 ;
        RECT -4.215 93.440 1.000 93.445 ;
        RECT 11.245 93.440 16.460 93.445 ;
        RECT 26.705 93.440 66.955 93.445 ;
        RECT -4.215 93.420 66.955 93.440 ;
        RECT 93.310 93.420 98.955 93.425 ;
        RECT 109.570 93.420 109.950 99.250 ;
        RECT 118.450 99.200 122.950 99.510 ;
        RECT 114.410 98.650 120.800 98.940 ;
        RECT 113.175 97.485 116.095 97.785 ;
        RECT 119.640 97.470 123.010 97.770 ;
        RECT 111.390 96.735 111.770 97.115 ;
        RECT 117.050 96.840 118.240 97.125 ;
        RECT 116.270 96.175 116.650 96.555 ;
        RECT 120.390 96.010 123.570 96.330 ;
        RECT 110.670 94.925 114.820 95.195 ;
        RECT 110.320 93.420 114.415 93.425 ;
        RECT -4.215 93.415 98.955 93.420 ;
        RECT 109.200 93.415 114.415 93.420 ;
        RECT -4.215 92.545 124.230 93.415 ;
        RECT 66.655 92.520 124.230 92.545 ;
        RECT 67.875 88.630 124.230 88.650 ;
        RECT -4.410 87.750 124.230 88.630 ;
        RECT -4.410 87.730 67.980 87.750 ;
        RECT -4.040 80.570 -3.660 87.730 ;
        RECT 1.535 83.275 1.915 83.655 ;
        RECT 8.435 83.265 8.815 83.645 ;
        RECT -1.140 82.850 0.600 83.140 ;
        RECT 5.360 82.770 7.970 83.195 ;
        RECT 7.545 80.330 10.650 80.605 ;
        RECT 11.420 80.570 11.800 87.730 ;
        RECT 64.860 86.745 93.635 86.765 ;
        RECT 28.060 86.480 93.635 86.745 ;
        RECT 28.060 86.460 65.610 86.480 ;
        RECT 95.305 86.460 102.010 86.760 ;
        RECT 31.765 85.550 32.965 85.930 ;
        RECT 34.720 85.335 36.995 85.845 ;
        RECT 39.620 85.335 41.920 85.845 ;
        RECT 44.215 85.335 46.495 85.845 ;
        RECT 51.290 85.650 52.525 86.030 ;
        RECT 68.165 85.570 69.620 85.950 ;
        RECT 73.315 85.355 75.590 85.865 ;
        RECT 78.215 85.355 80.515 85.865 ;
        RECT 82.810 85.355 85.090 85.865 ;
        RECT 91.860 85.670 93.140 86.050 ;
        RECT 52.705 85.295 53.085 85.330 ;
        RECT 91.300 85.315 91.680 85.350 ;
        RECT 31.205 85.190 31.585 85.230 ;
        RECT 31.135 84.885 33.970 85.190 ;
        RECT 49.950 84.985 53.085 85.295 ;
        RECT 69.800 85.210 70.180 85.250 ;
        RECT 52.705 84.950 53.085 84.985 ;
        RECT 69.730 84.905 72.565 85.210 ;
        RECT 88.545 85.005 91.680 85.315 ;
        RECT 91.300 84.970 91.680 85.005 ;
        RECT 31.205 84.850 31.585 84.885 ;
        RECT 69.800 84.870 70.180 84.905 ;
        RECT 13.250 83.475 16.655 83.915 ;
        RECT 16.995 83.275 17.375 83.655 ;
        RECT 19.710 83.315 20.090 83.695 ;
        RECT 23.895 83.265 24.275 83.645 ;
        RECT 31.765 83.250 35.025 83.630 ;
        RECT 35.765 83.250 39.025 83.630 ;
        RECT 45.265 83.250 48.525 83.630 ;
        RECT 49.265 83.250 52.525 83.630 ;
        RECT 68.325 83.270 69.620 83.650 ;
        RECT 74.360 83.270 77.620 83.650 ;
        RECT 78.360 83.270 79.545 83.650 ;
        RECT 81.810 83.270 83.120 83.650 ;
        RECT 83.860 83.270 87.120 83.650 ;
        RECT 91.860 83.270 92.875 83.650 ;
        RECT 95.940 83.515 99.355 83.935 ;
        RECT 99.685 83.295 100.065 83.675 ;
        RECT 102.400 83.335 102.780 83.715 ;
        RECT 106.585 83.285 106.965 83.665 ;
        RECT 14.320 82.850 16.060 83.140 ;
        RECT 18.110 82.800 19.310 83.090 ;
        RECT 20.820 82.770 23.415 83.145 ;
        RECT 25.030 82.865 25.410 83.245 ;
        RECT 31.205 82.550 31.585 82.930 ;
        RECT 35.205 82.550 35.585 82.930 ;
        RECT 39.205 82.885 39.585 82.930 ;
        RECT 44.705 82.885 45.085 82.930 ;
        RECT 39.155 82.570 45.090 82.885 ;
        RECT 39.205 82.550 39.585 82.570 ;
        RECT 44.705 82.550 45.085 82.570 ;
        RECT 48.705 82.550 49.085 82.930 ;
        RECT 52.705 82.550 53.085 82.930 ;
        RECT 69.800 82.570 70.180 82.950 ;
        RECT 73.800 82.570 74.180 82.950 ;
        RECT 77.800 82.905 78.180 82.950 ;
        RECT 83.300 82.905 83.680 82.950 ;
        RECT 77.750 82.590 83.685 82.905 ;
        RECT 77.800 82.570 78.180 82.590 ;
        RECT 83.300 82.570 83.680 82.590 ;
        RECT 87.300 82.570 87.680 82.950 ;
        RECT 91.300 82.570 91.680 82.950 ;
        RECT 97.010 82.870 98.750 83.160 ;
        RECT 100.800 82.820 102.000 83.110 ;
        RECT 103.510 82.780 106.140 83.235 ;
        RECT 107.720 82.885 108.100 83.265 ;
        RECT 61.890 81.945 82.665 82.320 ;
        RECT 32.430 81.335 59.740 81.675 ;
        RECT 12.045 80.630 19.305 80.930 ;
        RECT 12.600 80.095 16.685 80.365 ;
        RECT 23.005 80.330 26.755 80.605 ;
        RECT 60.920 80.590 92.885 80.980 ;
        RECT 105.695 80.350 108.825 80.625 ;
        RECT 109.570 80.590 109.950 87.750 ;
        RECT 110.810 85.290 117.550 85.590 ;
        RECT 111.400 83.495 114.855 83.935 ;
        RECT 117.860 83.335 118.240 83.715 ;
        RECT 116.260 82.820 117.460 83.110 ;
        RECT 123.180 82.885 123.560 83.265 ;
        RECT 110.215 82.110 126.135 82.410 ;
        RECT 110.750 81.365 127.695 81.665 ;
        RECT 57.765 80.225 85.325 80.235 ;
        RECT 28.060 80.205 46.730 80.215 ;
        RECT 57.765 80.205 94.330 80.225 ;
        RECT 28.060 79.915 94.330 80.205 ;
        RECT 28.060 79.895 58.080 79.915 ;
        RECT 111.945 79.455 116.075 79.755 ;
        RECT -4.040 73.605 -3.660 79.435 ;
        RECT 0.215 78.255 10.870 78.590 ;
        RECT 0.185 76.935 1.965 77.225 ;
        RECT 7.560 76.905 8.870 77.225 ;
        RECT -1.085 76.320 -0.705 76.700 ;
        RECT 5.370 76.350 5.750 76.730 ;
        RECT -3.290 73.605 0.805 73.610 ;
        RECT 11.420 73.605 11.800 79.435 ;
        RECT 62.985 79.225 94.730 79.245 ;
        RECT 16.260 78.835 22.650 79.125 ;
        RECT 27.530 78.975 94.730 79.225 ;
        RECT 27.530 78.955 63.440 78.975 ;
        RECT 98.950 78.855 105.340 79.145 ;
        RECT 15.675 78.255 26.180 78.590 ;
        RECT 51.150 78.390 61.700 78.725 ;
        RECT 98.365 78.275 108.845 78.610 ;
        RECT 31.745 77.750 35.045 78.130 ;
        RECT 35.745 77.750 39.045 78.130 ;
        RECT 45.245 77.750 48.545 78.130 ;
        RECT 49.245 77.750 52.545 78.130 ;
        RECT 68.335 77.770 69.640 78.150 ;
        RECT 74.340 77.770 77.640 78.150 ;
        RECT 78.340 77.770 79.700 78.150 ;
        RECT 81.675 77.770 83.140 78.150 ;
        RECT 83.840 77.770 87.140 78.150 ;
        RECT 91.840 77.770 93.020 78.150 ;
        RECT 31.205 77.405 31.585 77.440 ;
        RECT 13.240 76.920 13.620 77.300 ;
        RECT 15.645 76.935 17.425 77.225 ;
        RECT 18.900 77.025 20.090 77.310 ;
        RECT 23.020 76.905 24.330 77.225 ;
        RECT 30.940 77.095 33.950 77.405 ;
        RECT 31.205 77.060 31.585 77.095 ;
        RECT 35.205 77.060 36.295 77.440 ;
        RECT 39.205 77.435 39.585 77.440 ;
        RECT 36.725 77.070 39.590 77.435 ;
        RECT 44.705 77.415 45.085 77.440 ;
        RECT 44.690 77.095 46.835 77.415 ;
        RECT 39.205 77.060 39.585 77.070 ;
        RECT 44.705 77.060 45.085 77.095 ;
        RECT 47.750 77.060 49.085 77.440 ;
        RECT 52.705 77.420 53.085 77.440 ;
        RECT 69.800 77.425 70.180 77.460 ;
        RECT 50.240 77.100 53.150 77.420 ;
        RECT 69.535 77.115 72.545 77.425 ;
        RECT 52.705 77.060 53.085 77.100 ;
        RECT 69.800 77.080 70.180 77.115 ;
        RECT 73.800 77.080 74.890 77.460 ;
        RECT 77.800 77.455 78.180 77.460 ;
        RECT 75.320 77.090 78.185 77.455 ;
        RECT 83.300 77.435 83.680 77.460 ;
        RECT 83.285 77.115 85.430 77.435 ;
        RECT 77.800 77.080 78.180 77.090 ;
        RECT 83.300 77.080 83.680 77.115 ;
        RECT 86.345 77.080 87.680 77.460 ;
        RECT 91.300 77.440 91.680 77.460 ;
        RECT 88.835 77.120 91.745 77.440 ;
        RECT 91.300 77.080 91.680 77.120 ;
        RECT 95.930 76.940 96.310 77.320 ;
        RECT 98.335 76.955 100.115 77.245 ;
        RECT 101.590 77.045 102.780 77.330 ;
        RECT 105.710 76.925 107.020 77.245 ;
        RECT 14.375 76.320 14.755 76.700 ;
        RECT 18.120 76.360 18.500 76.740 ;
        RECT 20.830 76.350 21.210 76.730 ;
        RECT 22.240 76.195 25.420 76.515 ;
        RECT 97.065 76.340 97.445 76.720 ;
        RECT 100.810 76.380 101.190 76.760 ;
        RECT 103.520 76.370 103.900 76.750 ;
        RECT 104.930 76.215 108.110 76.535 ;
        RECT 31.745 75.750 33.030 76.130 ;
        RECT 51.060 75.750 52.545 76.130 ;
        RECT 68.150 75.770 69.640 76.150 ;
        RECT 91.840 75.770 92.915 76.150 ;
        RECT 31.205 75.060 32.295 75.440 ;
        RECT 33.250 75.070 34.770 75.430 ;
        RECT 35.690 75.065 48.540 75.400 ;
        RECT 52.705 75.395 53.085 75.440 ;
        RECT 51.970 75.095 53.280 75.395 ;
        RECT 52.705 75.060 53.085 75.095 ;
        RECT 69.800 75.080 70.890 75.460 ;
        RECT 71.845 75.090 73.365 75.450 ;
        RECT 74.285 75.085 87.135 75.420 ;
        RECT 91.300 75.415 91.680 75.460 ;
        RECT 90.565 75.115 91.875 75.415 ;
        RECT 91.300 75.080 91.680 75.115 ;
        RECT 60.360 74.550 93.310 74.585 ;
        RECT 28.060 74.220 93.310 74.550 ;
        RECT 28.060 74.200 61.140 74.220 ;
        RECT 95.105 74.210 99.365 74.565 ;
        RECT 93.310 73.625 98.955 73.630 ;
        RECT 109.570 73.625 109.950 79.455 ;
        RECT 118.450 79.405 122.950 79.715 ;
        RECT 114.410 78.855 120.800 79.145 ;
        RECT 113.175 77.690 116.095 77.990 ;
        RECT 119.640 77.675 123.010 77.975 ;
        RECT 111.390 76.940 111.770 77.320 ;
        RECT 117.050 77.045 118.240 77.330 ;
        RECT 116.270 76.380 116.650 76.760 ;
        RECT 120.390 76.215 123.570 76.535 ;
        RECT 110.670 75.130 114.820 75.400 ;
        RECT 110.320 73.625 114.415 73.630 ;
        RECT 66.655 73.620 98.955 73.625 ;
        RECT 109.200 73.620 114.415 73.625 ;
        RECT 12.170 73.605 16.265 73.610 ;
        RECT 66.655 73.605 124.230 73.620 ;
        RECT -4.410 73.600 0.805 73.605 ;
        RECT 11.050 73.600 16.265 73.605 ;
        RECT 26.510 73.600 124.230 73.605 ;
        RECT -4.410 72.725 124.230 73.600 ;
        RECT -4.410 72.705 66.760 72.725 ;
        RECT -4.540 68.895 67.850 68.920 ;
        RECT -4.540 68.020 124.150 68.895 ;
        RECT -4.170 60.860 -3.790 68.020 ;
        RECT 1.405 63.565 1.785 63.945 ;
        RECT 8.305 63.555 8.685 63.935 ;
        RECT -1.270 63.140 0.470 63.430 ;
        RECT 5.230 63.060 7.840 63.485 ;
        RECT 7.415 60.620 10.520 60.895 ;
        RECT 11.290 60.860 11.670 68.020 ;
        RECT 67.795 67.995 124.150 68.020 ;
        RECT 27.930 67.010 65.480 67.035 ;
        RECT 27.930 66.750 93.555 67.010 ;
        RECT 64.780 66.725 93.555 66.750 ;
        RECT 95.225 66.705 101.930 67.005 ;
        RECT 31.635 65.840 32.835 66.220 ;
        RECT 34.590 65.625 36.865 66.135 ;
        RECT 39.490 65.625 41.790 66.135 ;
        RECT 44.085 65.625 46.365 66.135 ;
        RECT 51.160 65.940 52.395 66.320 ;
        RECT 68.085 65.815 69.540 66.195 ;
        RECT 52.575 65.585 52.955 65.620 ;
        RECT 73.235 65.600 75.510 66.110 ;
        RECT 78.135 65.600 80.435 66.110 ;
        RECT 82.730 65.600 85.010 66.110 ;
        RECT 91.780 65.915 93.060 66.295 ;
        RECT 31.075 65.480 31.455 65.520 ;
        RECT 31.005 65.175 33.840 65.480 ;
        RECT 49.820 65.275 52.955 65.585 ;
        RECT 91.220 65.560 91.600 65.595 ;
        RECT 69.720 65.455 70.100 65.495 ;
        RECT 52.575 65.240 52.955 65.275 ;
        RECT 31.075 65.140 31.455 65.175 ;
        RECT 69.650 65.150 72.485 65.455 ;
        RECT 88.465 65.250 91.600 65.560 ;
        RECT 91.220 65.215 91.600 65.250 ;
        RECT 69.720 65.115 70.100 65.150 ;
        RECT 13.120 63.765 16.525 64.205 ;
        RECT 16.865 63.565 17.245 63.945 ;
        RECT 19.580 63.605 19.960 63.985 ;
        RECT 23.765 63.555 24.145 63.935 ;
        RECT 31.635 63.540 34.895 63.920 ;
        RECT 35.635 63.540 38.895 63.920 ;
        RECT 45.135 63.540 48.395 63.920 ;
        RECT 49.135 63.540 52.395 63.920 ;
        RECT 14.190 63.140 15.930 63.430 ;
        RECT 17.980 63.090 19.180 63.380 ;
        RECT 20.690 63.060 23.285 63.435 ;
        RECT 24.900 63.155 25.280 63.535 ;
        RECT 68.245 63.515 69.540 63.895 ;
        RECT 74.280 63.515 77.540 63.895 ;
        RECT 78.280 63.515 79.465 63.895 ;
        RECT 81.730 63.515 83.040 63.895 ;
        RECT 83.780 63.515 87.040 63.895 ;
        RECT 91.780 63.515 92.795 63.895 ;
        RECT 95.860 63.760 99.275 64.180 ;
        RECT 99.605 63.540 99.985 63.920 ;
        RECT 102.320 63.580 102.700 63.960 ;
        RECT 106.505 63.530 106.885 63.910 ;
        RECT 31.075 62.840 31.455 63.220 ;
        RECT 35.075 62.840 35.455 63.220 ;
        RECT 39.075 63.175 39.455 63.220 ;
        RECT 44.575 63.175 44.955 63.220 ;
        RECT 39.025 62.860 44.960 63.175 ;
        RECT 39.075 62.840 39.455 62.860 ;
        RECT 44.575 62.840 44.955 62.860 ;
        RECT 48.575 62.840 48.955 63.220 ;
        RECT 52.575 62.840 52.955 63.220 ;
        RECT 69.720 62.815 70.100 63.195 ;
        RECT 73.720 62.815 74.100 63.195 ;
        RECT 77.720 63.150 78.100 63.195 ;
        RECT 83.220 63.150 83.600 63.195 ;
        RECT 77.670 62.835 83.605 63.150 ;
        RECT 77.720 62.815 78.100 62.835 ;
        RECT 83.220 62.815 83.600 62.835 ;
        RECT 87.220 62.815 87.600 63.195 ;
        RECT 91.220 62.815 91.600 63.195 ;
        RECT 96.930 63.115 98.670 63.405 ;
        RECT 100.720 63.065 101.920 63.355 ;
        RECT 103.430 63.025 106.060 63.480 ;
        RECT 107.640 63.130 108.020 63.510 ;
        RECT 61.810 62.190 82.585 62.565 ;
        RECT 32.300 61.625 59.610 61.965 ;
        RECT 11.915 60.920 19.175 61.220 ;
        RECT 12.470 60.385 16.555 60.655 ;
        RECT 22.875 60.620 26.625 60.895 ;
        RECT 60.840 60.835 92.805 61.225 ;
        RECT 105.615 60.595 108.745 60.870 ;
        RECT 109.490 60.835 109.870 67.995 ;
        RECT 110.730 65.535 117.470 65.835 ;
        RECT 111.320 63.740 114.775 64.180 ;
        RECT 117.780 63.580 118.160 63.960 ;
        RECT 116.180 63.065 117.380 63.355 ;
        RECT 123.100 63.130 123.480 63.510 ;
        RECT 110.135 62.355 126.055 62.655 ;
        RECT 110.670 61.610 127.615 61.910 ;
        RECT 27.930 60.495 46.600 60.505 ;
        RECT 27.930 60.480 57.950 60.495 ;
        RECT 27.930 60.470 85.245 60.480 ;
        RECT 27.930 60.185 94.250 60.470 ;
        RECT 57.685 60.160 94.250 60.185 ;
        RECT -4.170 53.895 -3.790 59.725 ;
        RECT 0.085 58.545 10.740 58.880 ;
        RECT 0.055 57.225 1.835 57.515 ;
        RECT 7.430 57.195 8.740 57.515 ;
        RECT -1.215 56.610 -0.835 56.990 ;
        RECT 5.240 56.640 5.620 57.020 ;
        RECT -3.420 53.895 0.675 53.900 ;
        RECT 11.290 53.895 11.670 59.725 ;
        RECT 111.865 59.700 115.995 60.000 ;
        RECT 27.400 59.490 63.310 59.515 ;
        RECT 16.130 59.125 22.520 59.415 ;
        RECT 27.400 59.245 94.650 59.490 ;
        RECT 62.905 59.220 94.650 59.245 ;
        RECT 98.870 59.100 105.260 59.390 ;
        RECT 15.545 58.545 26.050 58.880 ;
        RECT 51.020 58.680 61.570 59.015 ;
        RECT 98.285 58.520 108.765 58.855 ;
        RECT 31.615 58.040 34.915 58.420 ;
        RECT 35.615 58.040 38.915 58.420 ;
        RECT 45.115 58.040 48.415 58.420 ;
        RECT 49.115 58.040 52.415 58.420 ;
        RECT 68.255 58.015 69.560 58.395 ;
        RECT 74.260 58.015 77.560 58.395 ;
        RECT 78.260 58.015 79.620 58.395 ;
        RECT 81.595 58.015 83.060 58.395 ;
        RECT 83.760 58.015 87.060 58.395 ;
        RECT 91.760 58.015 92.940 58.395 ;
        RECT 31.075 57.695 31.455 57.730 ;
        RECT 13.110 57.210 13.490 57.590 ;
        RECT 15.515 57.225 17.295 57.515 ;
        RECT 18.770 57.315 19.960 57.600 ;
        RECT 22.890 57.195 24.200 57.515 ;
        RECT 30.810 57.385 33.820 57.695 ;
        RECT 31.075 57.350 31.455 57.385 ;
        RECT 35.075 57.350 36.165 57.730 ;
        RECT 39.075 57.725 39.455 57.730 ;
        RECT 36.595 57.360 39.460 57.725 ;
        RECT 44.575 57.705 44.955 57.730 ;
        RECT 44.560 57.385 46.705 57.705 ;
        RECT 39.075 57.350 39.455 57.360 ;
        RECT 44.575 57.350 44.955 57.385 ;
        RECT 47.620 57.350 48.955 57.730 ;
        RECT 52.575 57.710 52.955 57.730 ;
        RECT 50.110 57.390 53.020 57.710 ;
        RECT 69.720 57.670 70.100 57.705 ;
        RECT 52.575 57.350 52.955 57.390 ;
        RECT 69.455 57.360 72.465 57.670 ;
        RECT 69.720 57.325 70.100 57.360 ;
        RECT 73.720 57.325 74.810 57.705 ;
        RECT 77.720 57.700 78.100 57.705 ;
        RECT 75.240 57.335 78.105 57.700 ;
        RECT 83.220 57.680 83.600 57.705 ;
        RECT 83.205 57.360 85.350 57.680 ;
        RECT 77.720 57.325 78.100 57.335 ;
        RECT 83.220 57.325 83.600 57.360 ;
        RECT 86.265 57.325 87.600 57.705 ;
        RECT 91.220 57.685 91.600 57.705 ;
        RECT 88.755 57.365 91.665 57.685 ;
        RECT 91.220 57.325 91.600 57.365 ;
        RECT 95.850 57.185 96.230 57.565 ;
        RECT 98.255 57.200 100.035 57.490 ;
        RECT 101.510 57.290 102.700 57.575 ;
        RECT 105.630 57.170 106.940 57.490 ;
        RECT 14.245 56.610 14.625 56.990 ;
        RECT 17.990 56.650 18.370 57.030 ;
        RECT 20.700 56.640 21.080 57.020 ;
        RECT 22.110 56.485 25.290 56.805 ;
        RECT 96.985 56.585 97.365 56.965 ;
        RECT 100.730 56.625 101.110 57.005 ;
        RECT 103.440 56.615 103.820 56.995 ;
        RECT 104.850 56.460 108.030 56.780 ;
        RECT 31.615 56.040 32.900 56.420 ;
        RECT 50.930 56.040 52.415 56.420 ;
        RECT 68.070 56.015 69.560 56.395 ;
        RECT 91.760 56.015 92.835 56.395 ;
        RECT 31.075 55.350 32.165 55.730 ;
        RECT 33.120 55.360 34.640 55.720 ;
        RECT 35.560 55.355 48.410 55.690 ;
        RECT 52.575 55.685 52.955 55.730 ;
        RECT 51.840 55.385 53.150 55.685 ;
        RECT 52.575 55.350 52.955 55.385 ;
        RECT 69.720 55.325 70.810 55.705 ;
        RECT 71.765 55.335 73.285 55.695 ;
        RECT 74.205 55.330 87.055 55.665 ;
        RECT 91.220 55.660 91.600 55.705 ;
        RECT 90.485 55.360 91.795 55.660 ;
        RECT 91.220 55.325 91.600 55.360 ;
        RECT 27.930 54.830 61.010 54.840 ;
        RECT 27.930 54.490 93.230 54.830 ;
        RECT 60.280 54.465 93.230 54.490 ;
        RECT 95.025 54.455 99.285 54.810 ;
        RECT 12.040 53.895 16.135 53.900 ;
        RECT -4.540 53.890 0.675 53.895 ;
        RECT 10.920 53.890 16.135 53.895 ;
        RECT 26.380 53.890 66.630 53.895 ;
        RECT -4.540 53.870 66.630 53.890 ;
        RECT 93.230 53.870 98.875 53.875 ;
        RECT 109.490 53.870 109.870 59.700 ;
        RECT 118.370 59.650 122.870 59.960 ;
        RECT 114.330 59.100 120.720 59.390 ;
        RECT 113.095 57.935 116.015 58.235 ;
        RECT 119.560 57.920 122.930 58.220 ;
        RECT 111.310 57.185 111.690 57.565 ;
        RECT 116.970 57.290 118.160 57.575 ;
        RECT 116.190 56.625 116.570 57.005 ;
        RECT 120.310 56.460 123.490 56.780 ;
        RECT 110.590 55.375 114.740 55.645 ;
        RECT 110.240 53.870 114.335 53.875 ;
        RECT -4.540 53.865 98.875 53.870 ;
        RECT 109.120 53.865 114.335 53.870 ;
        RECT -4.540 52.995 124.150 53.865 ;
        RECT 66.575 52.970 124.150 52.995 ;
        RECT 67.900 49.160 124.255 49.180 ;
        RECT -4.410 48.280 124.255 49.160 ;
        RECT -4.410 48.260 67.980 48.280 ;
        RECT -4.040 41.100 -3.660 48.260 ;
        RECT 1.535 43.805 1.915 44.185 ;
        RECT 8.435 43.795 8.815 44.175 ;
        RECT -1.140 43.380 0.600 43.670 ;
        RECT 5.360 43.300 7.970 43.725 ;
        RECT 7.545 40.860 10.650 41.135 ;
        RECT 11.420 41.100 11.800 48.260 ;
        RECT 64.885 47.275 93.660 47.295 ;
        RECT 28.060 47.010 93.660 47.275 ;
        RECT 28.060 46.990 65.610 47.010 ;
        RECT 95.330 46.990 102.035 47.290 ;
        RECT 31.765 46.080 32.965 46.460 ;
        RECT 34.720 45.865 36.995 46.375 ;
        RECT 39.620 45.865 41.920 46.375 ;
        RECT 44.215 45.865 46.495 46.375 ;
        RECT 51.290 46.180 52.525 46.560 ;
        RECT 68.190 46.100 69.645 46.480 ;
        RECT 73.340 45.885 75.615 46.395 ;
        RECT 78.240 45.885 80.540 46.395 ;
        RECT 82.835 45.885 85.115 46.395 ;
        RECT 91.885 46.200 93.165 46.580 ;
        RECT 52.705 45.825 53.085 45.860 ;
        RECT 91.325 45.845 91.705 45.880 ;
        RECT 31.205 45.720 31.585 45.760 ;
        RECT 31.135 45.415 33.970 45.720 ;
        RECT 49.950 45.515 53.085 45.825 ;
        RECT 69.825 45.740 70.205 45.780 ;
        RECT 52.705 45.480 53.085 45.515 ;
        RECT 69.755 45.435 72.590 45.740 ;
        RECT 88.570 45.535 91.705 45.845 ;
        RECT 91.325 45.500 91.705 45.535 ;
        RECT 31.205 45.380 31.585 45.415 ;
        RECT 69.825 45.400 70.205 45.435 ;
        RECT 13.250 44.005 16.655 44.445 ;
        RECT 16.995 43.805 17.375 44.185 ;
        RECT 19.710 43.845 20.090 44.225 ;
        RECT 23.895 43.795 24.275 44.175 ;
        RECT 31.765 43.780 35.025 44.160 ;
        RECT 35.765 43.780 39.025 44.160 ;
        RECT 45.265 43.780 48.525 44.160 ;
        RECT 49.265 43.780 52.525 44.160 ;
        RECT 68.350 43.800 69.645 44.180 ;
        RECT 74.385 43.800 77.645 44.180 ;
        RECT 78.385 43.800 79.570 44.180 ;
        RECT 81.835 43.800 83.145 44.180 ;
        RECT 83.885 43.800 87.145 44.180 ;
        RECT 91.885 43.800 92.900 44.180 ;
        RECT 95.965 44.045 99.380 44.465 ;
        RECT 99.710 43.825 100.090 44.205 ;
        RECT 102.425 43.865 102.805 44.245 ;
        RECT 106.610 43.815 106.990 44.195 ;
        RECT 14.320 43.380 16.060 43.670 ;
        RECT 18.110 43.330 19.310 43.620 ;
        RECT 20.820 43.300 23.415 43.675 ;
        RECT 25.030 43.395 25.410 43.775 ;
        RECT 31.205 43.080 31.585 43.460 ;
        RECT 35.205 43.080 35.585 43.460 ;
        RECT 39.205 43.415 39.585 43.460 ;
        RECT 44.705 43.415 45.085 43.460 ;
        RECT 39.155 43.100 45.090 43.415 ;
        RECT 39.205 43.080 39.585 43.100 ;
        RECT 44.705 43.080 45.085 43.100 ;
        RECT 48.705 43.080 49.085 43.460 ;
        RECT 52.705 43.080 53.085 43.460 ;
        RECT 69.825 43.100 70.205 43.480 ;
        RECT 73.825 43.100 74.205 43.480 ;
        RECT 77.825 43.435 78.205 43.480 ;
        RECT 83.325 43.435 83.705 43.480 ;
        RECT 77.775 43.120 83.710 43.435 ;
        RECT 77.825 43.100 78.205 43.120 ;
        RECT 83.325 43.100 83.705 43.120 ;
        RECT 87.325 43.100 87.705 43.480 ;
        RECT 91.325 43.100 91.705 43.480 ;
        RECT 97.035 43.400 98.775 43.690 ;
        RECT 100.825 43.350 102.025 43.640 ;
        RECT 103.535 43.310 106.165 43.765 ;
        RECT 107.745 43.415 108.125 43.795 ;
        RECT 61.915 42.475 82.690 42.850 ;
        RECT 32.430 41.865 59.740 42.205 ;
        RECT 12.045 41.160 19.305 41.460 ;
        RECT 12.600 40.625 16.685 40.895 ;
        RECT 23.005 40.860 26.755 41.135 ;
        RECT 60.945 41.120 92.910 41.510 ;
        RECT 105.720 40.880 108.850 41.155 ;
        RECT 109.595 41.120 109.975 48.280 ;
        RECT 110.835 45.820 117.575 46.120 ;
        RECT 111.425 44.025 114.880 44.465 ;
        RECT 117.885 43.865 118.265 44.245 ;
        RECT 116.285 43.350 117.485 43.640 ;
        RECT 123.205 43.415 123.585 43.795 ;
        RECT 110.240 42.640 126.160 42.940 ;
        RECT 110.775 41.895 127.720 42.195 ;
        RECT 57.790 40.755 85.350 40.765 ;
        RECT 28.060 40.735 46.730 40.745 ;
        RECT 57.790 40.735 94.355 40.755 ;
        RECT 28.060 40.445 94.355 40.735 ;
        RECT 28.060 40.425 58.080 40.445 ;
        RECT 111.970 39.985 116.100 40.285 ;
        RECT -4.040 34.135 -3.660 39.965 ;
        RECT 0.215 38.785 10.870 39.120 ;
        RECT 0.185 37.465 1.965 37.755 ;
        RECT 7.560 37.435 8.870 37.755 ;
        RECT -1.085 36.850 -0.705 37.230 ;
        RECT 5.370 36.880 5.750 37.260 ;
        RECT -3.290 34.135 0.805 34.140 ;
        RECT 11.420 34.135 11.800 39.965 ;
        RECT 63.010 39.755 94.755 39.775 ;
        RECT 16.260 39.365 22.650 39.655 ;
        RECT 27.530 39.505 94.755 39.755 ;
        RECT 27.530 39.485 63.440 39.505 ;
        RECT 98.975 39.385 105.365 39.675 ;
        RECT 15.675 38.785 26.180 39.120 ;
        RECT 51.150 38.920 61.700 39.255 ;
        RECT 98.390 38.805 108.870 39.140 ;
        RECT 31.745 38.280 35.045 38.660 ;
        RECT 35.745 38.280 39.045 38.660 ;
        RECT 45.245 38.280 48.545 38.660 ;
        RECT 49.245 38.280 52.545 38.660 ;
        RECT 68.360 38.300 69.665 38.680 ;
        RECT 74.365 38.300 77.665 38.680 ;
        RECT 78.365 38.300 79.725 38.680 ;
        RECT 81.700 38.300 83.165 38.680 ;
        RECT 83.865 38.300 87.165 38.680 ;
        RECT 91.865 38.300 93.045 38.680 ;
        RECT 31.205 37.935 31.585 37.970 ;
        RECT 13.240 37.450 13.620 37.830 ;
        RECT 15.645 37.465 17.425 37.755 ;
        RECT 18.900 37.555 20.090 37.840 ;
        RECT 23.020 37.435 24.330 37.755 ;
        RECT 30.940 37.625 33.950 37.935 ;
        RECT 31.205 37.590 31.585 37.625 ;
        RECT 35.205 37.590 36.295 37.970 ;
        RECT 39.205 37.965 39.585 37.970 ;
        RECT 36.725 37.600 39.590 37.965 ;
        RECT 44.705 37.945 45.085 37.970 ;
        RECT 44.690 37.625 46.835 37.945 ;
        RECT 39.205 37.590 39.585 37.600 ;
        RECT 44.705 37.590 45.085 37.625 ;
        RECT 47.750 37.590 49.085 37.970 ;
        RECT 52.705 37.950 53.085 37.970 ;
        RECT 69.825 37.955 70.205 37.990 ;
        RECT 50.240 37.630 53.150 37.950 ;
        RECT 69.560 37.645 72.570 37.955 ;
        RECT 52.705 37.590 53.085 37.630 ;
        RECT 69.825 37.610 70.205 37.645 ;
        RECT 73.825 37.610 74.915 37.990 ;
        RECT 77.825 37.985 78.205 37.990 ;
        RECT 75.345 37.620 78.210 37.985 ;
        RECT 83.325 37.965 83.705 37.990 ;
        RECT 83.310 37.645 85.455 37.965 ;
        RECT 77.825 37.610 78.205 37.620 ;
        RECT 83.325 37.610 83.705 37.645 ;
        RECT 86.370 37.610 87.705 37.990 ;
        RECT 91.325 37.970 91.705 37.990 ;
        RECT 88.860 37.650 91.770 37.970 ;
        RECT 91.325 37.610 91.705 37.650 ;
        RECT 95.955 37.470 96.335 37.850 ;
        RECT 98.360 37.485 100.140 37.775 ;
        RECT 101.615 37.575 102.805 37.860 ;
        RECT 105.735 37.455 107.045 37.775 ;
        RECT 14.375 36.850 14.755 37.230 ;
        RECT 18.120 36.890 18.500 37.270 ;
        RECT 20.830 36.880 21.210 37.260 ;
        RECT 22.240 36.725 25.420 37.045 ;
        RECT 97.090 36.870 97.470 37.250 ;
        RECT 100.835 36.910 101.215 37.290 ;
        RECT 103.545 36.900 103.925 37.280 ;
        RECT 104.955 36.745 108.135 37.065 ;
        RECT 31.745 36.280 33.030 36.660 ;
        RECT 51.060 36.280 52.545 36.660 ;
        RECT 68.175 36.300 69.665 36.680 ;
        RECT 91.865 36.300 92.940 36.680 ;
        RECT 31.205 35.590 32.295 35.970 ;
        RECT 33.250 35.600 34.770 35.960 ;
        RECT 35.690 35.595 48.540 35.930 ;
        RECT 52.705 35.925 53.085 35.970 ;
        RECT 51.970 35.625 53.280 35.925 ;
        RECT 52.705 35.590 53.085 35.625 ;
        RECT 69.825 35.610 70.915 35.990 ;
        RECT 71.870 35.620 73.390 35.980 ;
        RECT 74.310 35.615 87.160 35.950 ;
        RECT 91.325 35.945 91.705 35.990 ;
        RECT 90.590 35.645 91.900 35.945 ;
        RECT 91.325 35.610 91.705 35.645 ;
        RECT 60.385 35.080 93.335 35.115 ;
        RECT 28.060 34.750 93.335 35.080 ;
        RECT 28.060 34.730 61.140 34.750 ;
        RECT 95.130 34.740 99.390 35.095 ;
        RECT 93.335 34.155 98.980 34.160 ;
        RECT 109.595 34.155 109.975 39.985 ;
        RECT 118.475 39.935 122.975 40.245 ;
        RECT 114.435 39.385 120.825 39.675 ;
        RECT 113.200 38.220 116.120 38.520 ;
        RECT 119.665 38.205 123.035 38.505 ;
        RECT 111.415 37.470 111.795 37.850 ;
        RECT 117.075 37.575 118.265 37.860 ;
        RECT 116.295 36.910 116.675 37.290 ;
        RECT 120.415 36.745 123.595 37.065 ;
        RECT 110.695 35.660 114.845 35.930 ;
        RECT 110.345 34.155 114.440 34.160 ;
        RECT 66.680 34.150 98.980 34.155 ;
        RECT 109.225 34.150 114.440 34.155 ;
        RECT 12.170 34.135 16.265 34.140 ;
        RECT 66.680 34.135 124.255 34.150 ;
        RECT -4.410 34.130 0.805 34.135 ;
        RECT 11.050 34.130 16.265 34.135 ;
        RECT 26.510 34.130 124.255 34.135 ;
        RECT -4.410 33.255 124.255 34.130 ;
        RECT -4.410 33.235 66.760 33.255 ;
        RECT -4.460 29.210 67.930 29.350 ;
        RECT -4.460 28.450 124.255 29.210 ;
        RECT -4.090 21.290 -3.710 28.450 ;
        RECT 1.485 23.995 1.865 24.375 ;
        RECT 8.385 23.985 8.765 24.365 ;
        RECT -1.190 23.570 0.550 23.860 ;
        RECT 5.310 23.490 7.920 23.915 ;
        RECT 7.495 21.050 10.600 21.325 ;
        RECT 11.370 21.290 11.750 28.450 ;
        RECT 67.900 28.310 124.255 28.450 ;
        RECT 28.010 27.325 65.560 27.465 ;
        RECT 28.010 27.180 93.660 27.325 ;
        RECT 64.885 27.040 93.660 27.180 ;
        RECT 95.330 27.020 102.035 27.320 ;
        RECT 31.715 26.270 32.915 26.650 ;
        RECT 34.670 26.055 36.945 26.565 ;
        RECT 39.570 26.055 41.870 26.565 ;
        RECT 44.165 26.055 46.445 26.565 ;
        RECT 51.240 26.370 52.475 26.750 ;
        RECT 68.190 26.130 69.645 26.510 ;
        RECT 52.655 26.015 53.035 26.050 ;
        RECT 31.155 25.910 31.535 25.950 ;
        RECT 31.085 25.605 33.920 25.910 ;
        RECT 49.900 25.705 53.035 26.015 ;
        RECT 73.340 25.915 75.615 26.425 ;
        RECT 78.240 25.915 80.540 26.425 ;
        RECT 82.835 25.915 85.115 26.425 ;
        RECT 91.885 26.230 93.165 26.610 ;
        RECT 91.325 25.875 91.705 25.910 ;
        RECT 69.825 25.770 70.205 25.810 ;
        RECT 52.655 25.670 53.035 25.705 ;
        RECT 31.155 25.570 31.535 25.605 ;
        RECT 69.755 25.465 72.590 25.770 ;
        RECT 88.570 25.565 91.705 25.875 ;
        RECT 91.325 25.530 91.705 25.565 ;
        RECT 69.825 25.430 70.205 25.465 ;
        RECT 13.200 24.195 16.605 24.635 ;
        RECT 16.945 23.995 17.325 24.375 ;
        RECT 19.660 24.035 20.040 24.415 ;
        RECT 23.845 23.985 24.225 24.365 ;
        RECT 31.715 23.970 34.975 24.350 ;
        RECT 35.715 23.970 38.975 24.350 ;
        RECT 45.215 23.970 48.475 24.350 ;
        RECT 49.215 23.970 52.475 24.350 ;
        RECT 14.270 23.570 16.010 23.860 ;
        RECT 18.060 23.520 19.260 23.810 ;
        RECT 20.770 23.490 23.365 23.865 ;
        RECT 24.980 23.585 25.360 23.965 ;
        RECT 68.350 23.830 69.645 24.210 ;
        RECT 74.385 23.830 77.645 24.210 ;
        RECT 78.385 23.830 79.570 24.210 ;
        RECT 81.835 23.830 83.145 24.210 ;
        RECT 83.885 23.830 87.145 24.210 ;
        RECT 91.885 23.830 92.900 24.210 ;
        RECT 95.965 24.075 99.380 24.495 ;
        RECT 99.710 23.855 100.090 24.235 ;
        RECT 102.425 23.895 102.805 24.275 ;
        RECT 106.610 23.845 106.990 24.225 ;
        RECT 31.155 23.270 31.535 23.650 ;
        RECT 35.155 23.270 35.535 23.650 ;
        RECT 39.155 23.605 39.535 23.650 ;
        RECT 44.655 23.605 45.035 23.650 ;
        RECT 39.105 23.290 45.040 23.605 ;
        RECT 39.155 23.270 39.535 23.290 ;
        RECT 44.655 23.270 45.035 23.290 ;
        RECT 48.655 23.270 49.035 23.650 ;
        RECT 52.655 23.270 53.035 23.650 ;
        RECT 69.825 23.130 70.205 23.510 ;
        RECT 73.825 23.130 74.205 23.510 ;
        RECT 77.825 23.465 78.205 23.510 ;
        RECT 83.325 23.465 83.705 23.510 ;
        RECT 77.775 23.150 83.710 23.465 ;
        RECT 77.825 23.130 78.205 23.150 ;
        RECT 83.325 23.130 83.705 23.150 ;
        RECT 87.325 23.130 87.705 23.510 ;
        RECT 91.325 23.130 91.705 23.510 ;
        RECT 97.035 23.430 98.775 23.720 ;
        RECT 100.825 23.380 102.025 23.670 ;
        RECT 103.535 23.340 106.165 23.795 ;
        RECT 107.745 23.445 108.125 23.825 ;
        RECT 61.915 22.505 82.690 22.880 ;
        RECT 32.380 22.055 59.690 22.395 ;
        RECT 11.995 21.350 19.255 21.650 ;
        RECT 12.550 20.815 16.635 21.085 ;
        RECT 22.955 21.050 26.705 21.325 ;
        RECT 60.945 21.150 92.910 21.540 ;
        RECT 28.010 20.925 46.680 20.935 ;
        RECT 28.010 20.795 58.030 20.925 ;
        RECT 105.720 20.910 108.850 21.185 ;
        RECT 109.595 21.150 109.975 28.310 ;
        RECT 110.835 25.850 117.575 26.150 ;
        RECT 111.425 24.055 114.880 24.495 ;
        RECT 117.885 23.895 118.265 24.275 ;
        RECT 116.285 23.380 117.485 23.670 ;
        RECT 123.205 23.445 123.585 23.825 ;
        RECT 110.240 22.670 126.160 22.970 ;
        RECT 110.775 21.925 127.720 22.225 ;
        RECT 28.010 20.785 85.350 20.795 ;
        RECT 28.010 20.615 94.355 20.785 ;
        RECT 57.790 20.475 94.355 20.615 ;
        RECT -4.090 14.325 -3.710 20.155 ;
        RECT 0.165 18.975 10.820 19.310 ;
        RECT 0.135 17.655 1.915 17.945 ;
        RECT 7.510 17.625 8.820 17.945 ;
        RECT -1.135 17.040 -0.755 17.420 ;
        RECT 5.320 17.070 5.700 17.450 ;
        RECT -3.340 14.325 0.755 14.330 ;
        RECT 11.370 14.325 11.750 20.155 ;
        RECT 111.970 20.015 116.100 20.315 ;
        RECT 16.210 19.555 22.600 19.845 ;
        RECT 27.480 19.805 63.390 19.945 ;
        RECT 27.480 19.675 94.755 19.805 ;
        RECT 63.010 19.535 94.755 19.675 ;
        RECT 15.625 18.975 26.130 19.310 ;
        RECT 51.100 19.110 61.650 19.445 ;
        RECT 98.975 19.415 105.365 19.705 ;
        RECT 31.695 18.470 34.995 18.850 ;
        RECT 35.695 18.470 38.995 18.850 ;
        RECT 45.195 18.470 48.495 18.850 ;
        RECT 49.195 18.470 52.495 18.850 ;
        RECT 98.390 18.835 108.870 19.170 ;
        RECT 68.360 18.330 69.665 18.710 ;
        RECT 74.365 18.330 77.665 18.710 ;
        RECT 78.365 18.330 79.725 18.710 ;
        RECT 81.700 18.330 83.165 18.710 ;
        RECT 83.865 18.330 87.165 18.710 ;
        RECT 91.865 18.330 93.045 18.710 ;
        RECT 31.155 18.125 31.535 18.160 ;
        RECT 13.190 17.640 13.570 18.020 ;
        RECT 15.595 17.655 17.375 17.945 ;
        RECT 18.850 17.745 20.040 18.030 ;
        RECT 22.970 17.625 24.280 17.945 ;
        RECT 30.890 17.815 33.900 18.125 ;
        RECT 31.155 17.780 31.535 17.815 ;
        RECT 35.155 17.780 36.245 18.160 ;
        RECT 39.155 18.155 39.535 18.160 ;
        RECT 36.675 17.790 39.540 18.155 ;
        RECT 44.655 18.135 45.035 18.160 ;
        RECT 44.640 17.815 46.785 18.135 ;
        RECT 39.155 17.780 39.535 17.790 ;
        RECT 44.655 17.780 45.035 17.815 ;
        RECT 47.700 17.780 49.035 18.160 ;
        RECT 52.655 18.140 53.035 18.160 ;
        RECT 50.190 17.820 53.100 18.140 ;
        RECT 69.825 17.985 70.205 18.020 ;
        RECT 52.655 17.780 53.035 17.820 ;
        RECT 69.560 17.675 72.570 17.985 ;
        RECT 69.825 17.640 70.205 17.675 ;
        RECT 73.825 17.640 74.915 18.020 ;
        RECT 77.825 18.015 78.205 18.020 ;
        RECT 75.345 17.650 78.210 18.015 ;
        RECT 83.325 17.995 83.705 18.020 ;
        RECT 83.310 17.675 85.455 17.995 ;
        RECT 77.825 17.640 78.205 17.650 ;
        RECT 83.325 17.640 83.705 17.675 ;
        RECT 86.370 17.640 87.705 18.020 ;
        RECT 91.325 18.000 91.705 18.020 ;
        RECT 88.860 17.680 91.770 18.000 ;
        RECT 91.325 17.640 91.705 17.680 ;
        RECT 95.955 17.500 96.335 17.880 ;
        RECT 98.360 17.515 100.140 17.805 ;
        RECT 101.615 17.605 102.805 17.890 ;
        RECT 105.735 17.485 107.045 17.805 ;
        RECT 14.325 17.040 14.705 17.420 ;
        RECT 18.070 17.080 18.450 17.460 ;
        RECT 20.780 17.070 21.160 17.450 ;
        RECT 22.190 16.915 25.370 17.235 ;
        RECT 97.090 16.900 97.470 17.280 ;
        RECT 100.835 16.940 101.215 17.320 ;
        RECT 103.545 16.930 103.925 17.310 ;
        RECT 31.695 16.470 32.980 16.850 ;
        RECT 51.010 16.470 52.495 16.850 ;
        RECT 104.955 16.775 108.135 17.095 ;
        RECT 68.175 16.330 69.665 16.710 ;
        RECT 91.865 16.330 92.940 16.710 ;
        RECT 31.155 15.780 32.245 16.160 ;
        RECT 33.200 15.790 34.720 16.150 ;
        RECT 35.640 15.785 48.490 16.120 ;
        RECT 52.655 16.115 53.035 16.160 ;
        RECT 51.920 15.815 53.230 16.115 ;
        RECT 52.655 15.780 53.035 15.815 ;
        RECT 69.825 15.640 70.915 16.020 ;
        RECT 71.870 15.650 73.390 16.010 ;
        RECT 74.310 15.645 87.160 15.980 ;
        RECT 91.325 15.975 91.705 16.020 ;
        RECT 90.590 15.675 91.900 15.975 ;
        RECT 91.325 15.640 91.705 15.675 ;
        RECT 28.010 15.145 61.090 15.270 ;
        RECT 28.010 14.920 93.335 15.145 ;
        RECT 60.385 14.780 93.335 14.920 ;
        RECT 95.130 14.770 99.390 15.125 ;
        RECT 12.120 14.325 16.215 14.330 ;
        RECT -4.460 14.320 0.755 14.325 ;
        RECT 11.000 14.320 16.215 14.325 ;
        RECT 26.460 14.320 66.710 14.325 ;
        RECT -4.460 14.185 66.710 14.320 ;
        RECT 93.335 14.185 98.980 14.190 ;
        RECT 109.595 14.185 109.975 20.015 ;
        RECT 118.475 19.965 122.975 20.275 ;
        RECT 114.435 19.415 120.825 19.705 ;
        RECT 113.200 18.250 116.120 18.550 ;
        RECT 119.665 18.235 123.035 18.535 ;
        RECT 111.415 17.500 111.795 17.880 ;
        RECT 117.075 17.605 118.265 17.890 ;
        RECT 116.295 16.940 116.675 17.320 ;
        RECT 120.415 16.775 123.595 17.095 ;
        RECT 110.695 15.690 114.845 15.960 ;
        RECT 110.345 14.185 114.440 14.190 ;
        RECT -4.460 14.180 98.980 14.185 ;
        RECT 109.225 14.180 114.440 14.185 ;
        RECT -4.460 13.425 124.255 14.180 ;
        RECT 66.680 13.285 124.255 13.425 ;
        RECT -4.490 9.545 67.900 9.555 ;
        RECT -4.490 8.655 124.255 9.545 ;
        RECT -4.120 1.495 -3.740 8.655 ;
        RECT 1.455 4.200 1.835 4.580 ;
        RECT 8.355 4.190 8.735 4.570 ;
        RECT -1.220 3.775 0.520 4.065 ;
        RECT 5.280 3.695 7.890 4.120 ;
        RECT 7.465 1.255 10.570 1.530 ;
        RECT 11.340 1.495 11.720 8.655 ;
        RECT 67.900 8.645 124.255 8.655 ;
        RECT 27.980 7.660 65.530 7.670 ;
        RECT 27.980 7.385 93.660 7.660 ;
        RECT 64.885 7.375 93.660 7.385 ;
        RECT 95.330 7.355 102.035 7.655 ;
        RECT 31.685 6.475 32.885 6.855 ;
        RECT 34.640 6.260 36.915 6.770 ;
        RECT 39.540 6.260 41.840 6.770 ;
        RECT 44.135 6.260 46.415 6.770 ;
        RECT 51.210 6.575 52.445 6.955 ;
        RECT 68.190 6.465 69.645 6.845 ;
        RECT 52.625 6.220 53.005 6.255 ;
        RECT 73.340 6.250 75.615 6.760 ;
        RECT 78.240 6.250 80.540 6.760 ;
        RECT 82.835 6.250 85.115 6.760 ;
        RECT 91.885 6.565 93.165 6.945 ;
        RECT 31.125 6.115 31.505 6.155 ;
        RECT 31.055 5.810 33.890 6.115 ;
        RECT 49.870 5.910 53.005 6.220 ;
        RECT 91.325 6.210 91.705 6.245 ;
        RECT 69.825 6.105 70.205 6.145 ;
        RECT 52.625 5.875 53.005 5.910 ;
        RECT 31.125 5.775 31.505 5.810 ;
        RECT 69.755 5.800 72.590 6.105 ;
        RECT 88.570 5.900 91.705 6.210 ;
        RECT 91.325 5.865 91.705 5.900 ;
        RECT 69.825 5.765 70.205 5.800 ;
        RECT 13.170 4.400 16.575 4.840 ;
        RECT 16.915 4.200 17.295 4.580 ;
        RECT 19.630 4.240 20.010 4.620 ;
        RECT 23.815 4.190 24.195 4.570 ;
        RECT 31.685 4.175 34.945 4.555 ;
        RECT 35.685 4.175 38.945 4.555 ;
        RECT 45.185 4.175 48.445 4.555 ;
        RECT 49.185 4.175 52.445 4.555 ;
        RECT 14.240 3.775 15.980 4.065 ;
        RECT 18.030 3.725 19.230 4.015 ;
        RECT 20.740 3.695 23.335 4.070 ;
        RECT 24.950 3.790 25.330 4.170 ;
        RECT 68.350 4.165 69.645 4.545 ;
        RECT 74.385 4.165 77.645 4.545 ;
        RECT 78.385 4.165 79.570 4.545 ;
        RECT 81.835 4.165 83.145 4.545 ;
        RECT 83.885 4.165 87.145 4.545 ;
        RECT 91.885 4.165 92.900 4.545 ;
        RECT 95.965 4.410 99.380 4.830 ;
        RECT 99.710 4.190 100.090 4.570 ;
        RECT 102.425 4.230 102.805 4.610 ;
        RECT 106.610 4.180 106.990 4.560 ;
        RECT 31.125 3.475 31.505 3.855 ;
        RECT 35.125 3.475 35.505 3.855 ;
        RECT 39.125 3.810 39.505 3.855 ;
        RECT 44.625 3.810 45.005 3.855 ;
        RECT 39.075 3.495 45.010 3.810 ;
        RECT 39.125 3.475 39.505 3.495 ;
        RECT 44.625 3.475 45.005 3.495 ;
        RECT 48.625 3.475 49.005 3.855 ;
        RECT 52.625 3.475 53.005 3.855 ;
        RECT 69.825 3.465 70.205 3.845 ;
        RECT 73.825 3.465 74.205 3.845 ;
        RECT 77.825 3.800 78.205 3.845 ;
        RECT 83.325 3.800 83.705 3.845 ;
        RECT 77.775 3.485 83.710 3.800 ;
        RECT 77.825 3.465 78.205 3.485 ;
        RECT 83.325 3.465 83.705 3.485 ;
        RECT 87.325 3.465 87.705 3.845 ;
        RECT 91.325 3.465 91.705 3.845 ;
        RECT 97.035 3.765 98.775 4.055 ;
        RECT 100.825 3.715 102.025 4.005 ;
        RECT 103.535 3.675 106.165 4.130 ;
        RECT 107.745 3.780 108.125 4.160 ;
        RECT 61.915 2.840 82.690 3.215 ;
        RECT 32.350 2.260 59.660 2.600 ;
        RECT 11.965 1.555 19.225 1.855 ;
        RECT 12.520 1.020 16.605 1.290 ;
        RECT 22.925 1.255 26.675 1.530 ;
        RECT 60.945 1.485 92.910 1.875 ;
        RECT 105.720 1.245 108.850 1.520 ;
        RECT 109.595 1.485 109.975 8.645 ;
        RECT 110.835 6.185 117.575 6.485 ;
        RECT 111.425 4.390 114.880 4.830 ;
        RECT 117.885 4.230 118.265 4.610 ;
        RECT 116.285 3.715 117.485 4.005 ;
        RECT 123.205 3.780 123.585 4.160 ;
        RECT 110.240 3.005 126.160 3.305 ;
        RECT 110.775 2.260 127.720 2.560 ;
        RECT 27.980 1.130 46.650 1.140 ;
        RECT 27.980 1.120 85.350 1.130 ;
        RECT 27.980 0.820 94.355 1.120 ;
        RECT 57.790 0.810 94.355 0.820 ;
        RECT -4.120 -5.470 -3.740 0.360 ;
        RECT 0.135 -0.820 10.790 -0.485 ;
        RECT 0.105 -2.140 1.885 -1.850 ;
        RECT 7.480 -2.170 8.790 -1.850 ;
        RECT -1.165 -2.755 -0.785 -2.375 ;
        RECT 5.290 -2.725 5.670 -2.345 ;
        RECT -3.370 -5.470 0.725 -5.465 ;
        RECT 11.340 -5.470 11.720 0.360 ;
        RECT 111.970 0.350 116.100 0.650 ;
        RECT 27.450 0.140 63.360 0.150 ;
        RECT 16.180 -0.240 22.570 0.050 ;
        RECT 27.450 -0.120 94.755 0.140 ;
        RECT 63.010 -0.130 94.755 -0.120 ;
        RECT 98.975 -0.250 105.365 0.040 ;
        RECT 15.595 -0.820 26.100 -0.485 ;
        RECT 51.070 -0.685 61.620 -0.350 ;
        RECT 98.390 -0.830 108.870 -0.495 ;
        RECT 31.665 -1.325 34.965 -0.945 ;
        RECT 35.665 -1.325 38.965 -0.945 ;
        RECT 45.165 -1.325 48.465 -0.945 ;
        RECT 49.165 -1.325 52.465 -0.945 ;
        RECT 68.360 -1.335 69.665 -0.955 ;
        RECT 74.365 -1.335 77.665 -0.955 ;
        RECT 78.365 -1.335 79.725 -0.955 ;
        RECT 81.700 -1.335 83.165 -0.955 ;
        RECT 83.865 -1.335 87.165 -0.955 ;
        RECT 91.865 -1.335 93.045 -0.955 ;
        RECT 31.125 -1.670 31.505 -1.635 ;
        RECT 13.160 -2.155 13.540 -1.775 ;
        RECT 15.565 -2.140 17.345 -1.850 ;
        RECT 18.820 -2.050 20.010 -1.765 ;
        RECT 22.940 -2.170 24.250 -1.850 ;
        RECT 30.860 -1.980 33.870 -1.670 ;
        RECT 31.125 -2.015 31.505 -1.980 ;
        RECT 35.125 -2.015 36.215 -1.635 ;
        RECT 39.125 -1.640 39.505 -1.635 ;
        RECT 36.645 -2.005 39.510 -1.640 ;
        RECT 44.625 -1.660 45.005 -1.635 ;
        RECT 44.610 -1.980 46.755 -1.660 ;
        RECT 39.125 -2.015 39.505 -2.005 ;
        RECT 44.625 -2.015 45.005 -1.980 ;
        RECT 47.670 -2.015 49.005 -1.635 ;
        RECT 52.625 -1.655 53.005 -1.635 ;
        RECT 50.160 -1.975 53.070 -1.655 ;
        RECT 69.825 -1.680 70.205 -1.645 ;
        RECT 52.625 -2.015 53.005 -1.975 ;
        RECT 69.560 -1.990 72.570 -1.680 ;
        RECT 69.825 -2.025 70.205 -1.990 ;
        RECT 73.825 -2.025 74.915 -1.645 ;
        RECT 77.825 -1.650 78.205 -1.645 ;
        RECT 75.345 -2.015 78.210 -1.650 ;
        RECT 83.325 -1.670 83.705 -1.645 ;
        RECT 83.310 -1.990 85.455 -1.670 ;
        RECT 77.825 -2.025 78.205 -2.015 ;
        RECT 83.325 -2.025 83.705 -1.990 ;
        RECT 86.370 -2.025 87.705 -1.645 ;
        RECT 91.325 -1.665 91.705 -1.645 ;
        RECT 88.860 -1.985 91.770 -1.665 ;
        RECT 91.325 -2.025 91.705 -1.985 ;
        RECT 95.955 -2.165 96.335 -1.785 ;
        RECT 98.360 -2.150 100.140 -1.860 ;
        RECT 101.615 -2.060 102.805 -1.775 ;
        RECT 105.735 -2.180 107.045 -1.860 ;
        RECT 14.295 -2.755 14.675 -2.375 ;
        RECT 18.040 -2.715 18.420 -2.335 ;
        RECT 20.750 -2.725 21.130 -2.345 ;
        RECT 22.160 -2.880 25.340 -2.560 ;
        RECT 97.090 -2.765 97.470 -2.385 ;
        RECT 100.835 -2.725 101.215 -2.345 ;
        RECT 103.545 -2.735 103.925 -2.355 ;
        RECT 104.955 -2.890 108.135 -2.570 ;
        RECT 31.665 -3.325 32.950 -2.945 ;
        RECT 50.980 -3.325 52.465 -2.945 ;
        RECT 68.175 -3.335 69.665 -2.955 ;
        RECT 91.865 -3.335 92.940 -2.955 ;
        RECT 31.125 -4.015 32.215 -3.635 ;
        RECT 33.170 -4.005 34.690 -3.645 ;
        RECT 35.610 -4.010 48.460 -3.675 ;
        RECT 52.625 -3.680 53.005 -3.635 ;
        RECT 51.890 -3.980 53.200 -3.680 ;
        RECT 52.625 -4.015 53.005 -3.980 ;
        RECT 69.825 -4.025 70.915 -3.645 ;
        RECT 71.870 -4.015 73.390 -3.655 ;
        RECT 74.310 -4.020 87.160 -3.685 ;
        RECT 91.325 -3.690 91.705 -3.645 ;
        RECT 90.590 -3.990 91.900 -3.690 ;
        RECT 91.325 -4.025 91.705 -3.990 ;
        RECT 60.385 -4.525 93.335 -4.520 ;
        RECT 27.980 -4.875 93.335 -4.525 ;
        RECT 60.385 -4.885 93.335 -4.875 ;
        RECT 95.130 -4.895 99.390 -4.540 ;
        RECT 12.090 -5.470 16.185 -5.465 ;
        RECT -4.490 -5.475 0.725 -5.470 ;
        RECT 10.970 -5.475 16.185 -5.470 ;
        RECT 26.430 -5.475 66.680 -5.470 ;
        RECT -4.490 -5.480 66.680 -5.475 ;
        RECT 93.335 -5.480 98.980 -5.475 ;
        RECT 109.595 -5.480 109.975 0.350 ;
        RECT 118.475 0.300 122.975 0.610 ;
        RECT 114.435 -0.250 120.825 0.040 ;
        RECT 113.200 -1.415 116.120 -1.115 ;
        RECT 119.665 -1.430 123.035 -1.130 ;
        RECT 111.415 -2.165 111.795 -1.785 ;
        RECT 117.075 -2.060 118.265 -1.775 ;
        RECT 116.295 -2.725 116.675 -2.345 ;
        RECT 120.415 -2.890 123.595 -2.570 ;
        RECT 110.695 -3.975 114.845 -3.705 ;
        RECT 110.345 -5.480 114.440 -5.475 ;
        RECT -4.490 -5.485 98.980 -5.480 ;
        RECT 109.225 -5.485 114.440 -5.480 ;
        RECT -4.490 -6.370 124.255 -5.485 ;
        RECT 66.680 -6.380 124.255 -6.370 ;
        RECT -4.340 -10.295 68.050 -10.240 ;
        RECT -4.340 -11.140 124.295 -10.295 ;
        RECT -3.970 -18.300 -3.590 -11.140 ;
        RECT 1.605 -15.595 1.985 -15.215 ;
        RECT 8.505 -15.605 8.885 -15.225 ;
        RECT -1.070 -16.020 0.670 -15.730 ;
        RECT 5.430 -16.100 8.040 -15.675 ;
        RECT 7.615 -18.540 10.720 -18.265 ;
        RECT 11.490 -18.300 11.870 -11.140 ;
        RECT 67.940 -11.195 124.295 -11.140 ;
        RECT 28.130 -12.180 65.680 -12.125 ;
        RECT 28.130 -12.410 93.700 -12.180 ;
        RECT 64.925 -12.465 93.700 -12.410 ;
        RECT 95.370 -12.485 102.075 -12.185 ;
        RECT 31.835 -13.320 33.035 -12.940 ;
        RECT 34.790 -13.535 37.065 -13.025 ;
        RECT 39.690 -13.535 41.990 -13.025 ;
        RECT 44.285 -13.535 46.565 -13.025 ;
        RECT 51.360 -13.220 52.595 -12.840 ;
        RECT 68.230 -13.375 69.685 -12.995 ;
        RECT 52.775 -13.575 53.155 -13.540 ;
        RECT 31.275 -13.680 31.655 -13.640 ;
        RECT 31.205 -13.985 34.040 -13.680 ;
        RECT 50.020 -13.885 53.155 -13.575 ;
        RECT 73.380 -13.590 75.655 -13.080 ;
        RECT 78.280 -13.590 80.580 -13.080 ;
        RECT 82.875 -13.590 85.155 -13.080 ;
        RECT 91.925 -13.275 93.205 -12.895 ;
        RECT 91.365 -13.630 91.745 -13.595 ;
        RECT 69.865 -13.735 70.245 -13.695 ;
        RECT 52.775 -13.920 53.155 -13.885 ;
        RECT 31.275 -14.020 31.655 -13.985 ;
        RECT 69.795 -14.040 72.630 -13.735 ;
        RECT 88.610 -13.940 91.745 -13.630 ;
        RECT 91.365 -13.975 91.745 -13.940 ;
        RECT 69.865 -14.075 70.245 -14.040 ;
        RECT 13.320 -15.395 16.725 -14.955 ;
        RECT 17.065 -15.595 17.445 -15.215 ;
        RECT 19.780 -15.555 20.160 -15.175 ;
        RECT 23.965 -15.605 24.345 -15.225 ;
        RECT 31.835 -15.620 35.095 -15.240 ;
        RECT 35.835 -15.620 39.095 -15.240 ;
        RECT 45.335 -15.620 48.595 -15.240 ;
        RECT 49.335 -15.620 52.595 -15.240 ;
        RECT 14.390 -16.020 16.130 -15.730 ;
        RECT 18.180 -16.070 19.380 -15.780 ;
        RECT 20.890 -16.100 23.485 -15.725 ;
        RECT 25.100 -16.005 25.480 -15.625 ;
        RECT 68.390 -15.675 69.685 -15.295 ;
        RECT 74.425 -15.675 77.685 -15.295 ;
        RECT 78.425 -15.675 79.610 -15.295 ;
        RECT 81.875 -15.675 83.185 -15.295 ;
        RECT 83.925 -15.675 87.185 -15.295 ;
        RECT 91.925 -15.675 92.940 -15.295 ;
        RECT 96.005 -15.430 99.420 -15.010 ;
        RECT 99.750 -15.650 100.130 -15.270 ;
        RECT 102.465 -15.610 102.845 -15.230 ;
        RECT 106.650 -15.660 107.030 -15.280 ;
        RECT 31.275 -16.320 31.655 -15.940 ;
        RECT 35.275 -16.320 35.655 -15.940 ;
        RECT 39.275 -15.985 39.655 -15.940 ;
        RECT 44.775 -15.985 45.155 -15.940 ;
        RECT 39.225 -16.300 45.160 -15.985 ;
        RECT 39.275 -16.320 39.655 -16.300 ;
        RECT 44.775 -16.320 45.155 -16.300 ;
        RECT 48.775 -16.320 49.155 -15.940 ;
        RECT 52.775 -16.320 53.155 -15.940 ;
        RECT 69.865 -16.375 70.245 -15.995 ;
        RECT 73.865 -16.375 74.245 -15.995 ;
        RECT 77.865 -16.040 78.245 -15.995 ;
        RECT 83.365 -16.040 83.745 -15.995 ;
        RECT 77.815 -16.355 83.750 -16.040 ;
        RECT 77.865 -16.375 78.245 -16.355 ;
        RECT 83.365 -16.375 83.745 -16.355 ;
        RECT 87.365 -16.375 87.745 -15.995 ;
        RECT 91.365 -16.375 91.745 -15.995 ;
        RECT 97.075 -16.075 98.815 -15.785 ;
        RECT 100.865 -16.125 102.065 -15.835 ;
        RECT 103.575 -16.165 106.205 -15.710 ;
        RECT 107.785 -16.060 108.165 -15.680 ;
        RECT 61.955 -17.000 82.730 -16.625 ;
        RECT 32.500 -17.535 59.810 -17.195 ;
        RECT 12.115 -18.240 19.375 -17.940 ;
        RECT 12.670 -18.775 16.755 -18.505 ;
        RECT 23.075 -18.540 26.825 -18.265 ;
        RECT 60.985 -18.355 92.950 -17.965 ;
        RECT 105.760 -18.595 108.890 -18.320 ;
        RECT 109.635 -18.355 110.015 -11.195 ;
        RECT 110.875 -13.655 117.615 -13.355 ;
        RECT 111.465 -15.450 114.920 -15.010 ;
        RECT 117.925 -15.610 118.305 -15.230 ;
        RECT 116.325 -16.125 117.525 -15.835 ;
        RECT 123.245 -16.060 123.625 -15.680 ;
        RECT 110.280 -16.835 126.200 -16.535 ;
        RECT 110.815 -17.580 127.760 -17.280 ;
        RECT 28.130 -18.665 46.800 -18.655 ;
        RECT 28.130 -18.710 58.150 -18.665 ;
        RECT 28.130 -18.720 85.390 -18.710 ;
        RECT 28.130 -18.975 94.395 -18.720 ;
        RECT 57.830 -19.030 94.395 -18.975 ;
        RECT -3.970 -25.265 -3.590 -19.435 ;
        RECT 0.285 -20.615 10.940 -20.280 ;
        RECT 0.255 -21.935 2.035 -21.645 ;
        RECT 7.630 -21.965 8.940 -21.645 ;
        RECT -1.015 -22.550 -0.635 -22.170 ;
        RECT 5.440 -22.520 5.820 -22.140 ;
        RECT -3.220 -25.265 0.875 -25.260 ;
        RECT 11.490 -25.265 11.870 -19.435 ;
        RECT 112.010 -19.490 116.140 -19.190 ;
        RECT 27.600 -19.700 63.510 -19.645 ;
        RECT 16.330 -20.035 22.720 -19.745 ;
        RECT 27.600 -19.915 94.795 -19.700 ;
        RECT 63.050 -19.970 94.795 -19.915 ;
        RECT 99.015 -20.090 105.405 -19.800 ;
        RECT 15.745 -20.615 26.250 -20.280 ;
        RECT 51.220 -20.480 61.770 -20.145 ;
        RECT 98.430 -20.670 108.910 -20.335 ;
        RECT 31.815 -21.120 35.115 -20.740 ;
        RECT 35.815 -21.120 39.115 -20.740 ;
        RECT 45.315 -21.120 48.615 -20.740 ;
        RECT 49.315 -21.120 52.615 -20.740 ;
        RECT 68.400 -21.175 69.705 -20.795 ;
        RECT 74.405 -21.175 77.705 -20.795 ;
        RECT 78.405 -21.175 79.765 -20.795 ;
        RECT 81.740 -21.175 83.205 -20.795 ;
        RECT 83.905 -21.175 87.205 -20.795 ;
        RECT 91.905 -21.175 93.085 -20.795 ;
        RECT 31.275 -21.465 31.655 -21.430 ;
        RECT 13.310 -21.950 13.690 -21.570 ;
        RECT 15.715 -21.935 17.495 -21.645 ;
        RECT 18.970 -21.845 20.160 -21.560 ;
        RECT 23.090 -21.965 24.400 -21.645 ;
        RECT 31.010 -21.775 34.020 -21.465 ;
        RECT 31.275 -21.810 31.655 -21.775 ;
        RECT 35.275 -21.810 36.365 -21.430 ;
        RECT 39.275 -21.435 39.655 -21.430 ;
        RECT 36.795 -21.800 39.660 -21.435 ;
        RECT 44.775 -21.455 45.155 -21.430 ;
        RECT 44.760 -21.775 46.905 -21.455 ;
        RECT 39.275 -21.810 39.655 -21.800 ;
        RECT 44.775 -21.810 45.155 -21.775 ;
        RECT 47.820 -21.810 49.155 -21.430 ;
        RECT 52.775 -21.450 53.155 -21.430 ;
        RECT 50.310 -21.770 53.220 -21.450 ;
        RECT 69.865 -21.520 70.245 -21.485 ;
        RECT 52.775 -21.810 53.155 -21.770 ;
        RECT 69.600 -21.830 72.610 -21.520 ;
        RECT 69.865 -21.865 70.245 -21.830 ;
        RECT 73.865 -21.865 74.955 -21.485 ;
        RECT 77.865 -21.490 78.245 -21.485 ;
        RECT 75.385 -21.855 78.250 -21.490 ;
        RECT 83.365 -21.510 83.745 -21.485 ;
        RECT 83.350 -21.830 85.495 -21.510 ;
        RECT 77.865 -21.865 78.245 -21.855 ;
        RECT 83.365 -21.865 83.745 -21.830 ;
        RECT 86.410 -21.865 87.745 -21.485 ;
        RECT 91.365 -21.505 91.745 -21.485 ;
        RECT 88.900 -21.825 91.810 -21.505 ;
        RECT 91.365 -21.865 91.745 -21.825 ;
        RECT 95.995 -22.005 96.375 -21.625 ;
        RECT 98.400 -21.990 100.180 -21.700 ;
        RECT 101.655 -21.900 102.845 -21.615 ;
        RECT 105.775 -22.020 107.085 -21.700 ;
        RECT 14.445 -22.550 14.825 -22.170 ;
        RECT 18.190 -22.510 18.570 -22.130 ;
        RECT 20.900 -22.520 21.280 -22.140 ;
        RECT 22.310 -22.675 25.490 -22.355 ;
        RECT 97.130 -22.605 97.510 -22.225 ;
        RECT 100.875 -22.565 101.255 -22.185 ;
        RECT 103.585 -22.575 103.965 -22.195 ;
        RECT 104.995 -22.730 108.175 -22.410 ;
        RECT 31.815 -23.120 33.100 -22.740 ;
        RECT 51.130 -23.120 52.615 -22.740 ;
        RECT 68.215 -23.175 69.705 -22.795 ;
        RECT 91.905 -23.175 92.980 -22.795 ;
        RECT 31.275 -23.810 32.365 -23.430 ;
        RECT 33.320 -23.800 34.840 -23.440 ;
        RECT 35.760 -23.805 48.610 -23.470 ;
        RECT 52.775 -23.475 53.155 -23.430 ;
        RECT 52.040 -23.775 53.350 -23.475 ;
        RECT 52.775 -23.810 53.155 -23.775 ;
        RECT 69.865 -23.865 70.955 -23.485 ;
        RECT 71.910 -23.855 73.430 -23.495 ;
        RECT 74.350 -23.860 87.200 -23.525 ;
        RECT 91.365 -23.530 91.745 -23.485 ;
        RECT 90.630 -23.830 91.940 -23.530 ;
        RECT 91.365 -23.865 91.745 -23.830 ;
        RECT 28.130 -24.360 61.210 -24.320 ;
        RECT 28.130 -24.670 93.375 -24.360 ;
        RECT 60.425 -24.725 93.375 -24.670 ;
        RECT 95.170 -24.735 99.430 -24.380 ;
        RECT 12.240 -25.265 16.335 -25.260 ;
        RECT -4.340 -25.270 0.875 -25.265 ;
        RECT 11.120 -25.270 16.335 -25.265 ;
        RECT 26.580 -25.270 66.830 -25.265 ;
        RECT -4.340 -25.320 66.830 -25.270 ;
        RECT 93.375 -25.320 99.020 -25.315 ;
        RECT 109.635 -25.320 110.015 -19.490 ;
        RECT 118.515 -19.540 123.015 -19.230 ;
        RECT 114.475 -20.090 120.865 -19.800 ;
        RECT 113.240 -21.255 116.160 -20.955 ;
        RECT 119.705 -21.270 123.075 -20.970 ;
        RECT 111.455 -22.005 111.835 -21.625 ;
        RECT 117.115 -21.900 118.305 -21.615 ;
        RECT 116.335 -22.565 116.715 -22.185 ;
        RECT 120.455 -22.730 123.635 -22.410 ;
        RECT 110.735 -23.815 114.885 -23.545 ;
        RECT 110.385 -25.320 114.480 -25.315 ;
        RECT -4.340 -25.325 99.020 -25.320 ;
        RECT 109.265 -25.325 114.480 -25.320 ;
        RECT -4.340 -26.165 124.295 -25.325 ;
        RECT 66.720 -26.220 124.295 -26.165 ;
        RECT -4.385 -30.020 68.005 -29.930 ;
        RECT -4.385 -30.830 124.095 -30.020 ;
        RECT -4.015 -37.990 -3.635 -30.830 ;
        RECT 1.560 -35.285 1.940 -34.905 ;
        RECT 8.460 -35.295 8.840 -34.915 ;
        RECT -1.115 -35.710 0.625 -35.420 ;
        RECT 5.385 -35.790 7.995 -35.365 ;
        RECT 7.570 -38.230 10.675 -37.955 ;
        RECT 11.445 -37.990 11.825 -30.830 ;
        RECT 67.740 -30.920 124.095 -30.830 ;
        RECT 28.085 -31.905 65.635 -31.815 ;
        RECT 28.085 -32.100 93.500 -31.905 ;
        RECT 64.725 -32.190 93.500 -32.100 ;
        RECT 95.170 -32.210 101.875 -31.910 ;
        RECT 31.790 -33.010 32.990 -32.630 ;
        RECT 34.745 -33.225 37.020 -32.715 ;
        RECT 39.645 -33.225 41.945 -32.715 ;
        RECT 44.240 -33.225 46.520 -32.715 ;
        RECT 51.315 -32.910 52.550 -32.530 ;
        RECT 68.030 -33.100 69.485 -32.720 ;
        RECT 52.730 -33.265 53.110 -33.230 ;
        RECT 31.230 -33.370 31.610 -33.330 ;
        RECT 31.160 -33.675 33.995 -33.370 ;
        RECT 49.975 -33.575 53.110 -33.265 ;
        RECT 73.180 -33.315 75.455 -32.805 ;
        RECT 78.080 -33.315 80.380 -32.805 ;
        RECT 82.675 -33.315 84.955 -32.805 ;
        RECT 91.725 -33.000 93.005 -32.620 ;
        RECT 91.165 -33.355 91.545 -33.320 ;
        RECT 69.665 -33.460 70.045 -33.420 ;
        RECT 52.730 -33.610 53.110 -33.575 ;
        RECT 31.230 -33.710 31.610 -33.675 ;
        RECT 69.595 -33.765 72.430 -33.460 ;
        RECT 88.410 -33.665 91.545 -33.355 ;
        RECT 91.165 -33.700 91.545 -33.665 ;
        RECT 69.665 -33.800 70.045 -33.765 ;
        RECT 13.275 -35.085 16.680 -34.645 ;
        RECT 17.020 -35.285 17.400 -34.905 ;
        RECT 19.735 -35.245 20.115 -34.865 ;
        RECT 23.920 -35.295 24.300 -34.915 ;
        RECT 31.790 -35.310 35.050 -34.930 ;
        RECT 35.790 -35.310 39.050 -34.930 ;
        RECT 45.290 -35.310 48.550 -34.930 ;
        RECT 49.290 -35.310 52.550 -34.930 ;
        RECT 14.345 -35.710 16.085 -35.420 ;
        RECT 18.135 -35.760 19.335 -35.470 ;
        RECT 20.845 -35.790 23.440 -35.415 ;
        RECT 25.055 -35.695 25.435 -35.315 ;
        RECT 68.190 -35.400 69.485 -35.020 ;
        RECT 74.225 -35.400 77.485 -35.020 ;
        RECT 78.225 -35.400 79.410 -35.020 ;
        RECT 81.675 -35.400 82.985 -35.020 ;
        RECT 83.725 -35.400 86.985 -35.020 ;
        RECT 91.725 -35.400 92.740 -35.020 ;
        RECT 95.805 -35.155 99.220 -34.735 ;
        RECT 99.550 -35.375 99.930 -34.995 ;
        RECT 102.265 -35.335 102.645 -34.955 ;
        RECT 106.450 -35.385 106.830 -35.005 ;
        RECT 31.230 -36.010 31.610 -35.630 ;
        RECT 35.230 -36.010 35.610 -35.630 ;
        RECT 39.230 -35.675 39.610 -35.630 ;
        RECT 44.730 -35.675 45.110 -35.630 ;
        RECT 39.180 -35.990 45.115 -35.675 ;
        RECT 39.230 -36.010 39.610 -35.990 ;
        RECT 44.730 -36.010 45.110 -35.990 ;
        RECT 48.730 -36.010 49.110 -35.630 ;
        RECT 52.730 -36.010 53.110 -35.630 ;
        RECT 69.665 -36.100 70.045 -35.720 ;
        RECT 73.665 -36.100 74.045 -35.720 ;
        RECT 77.665 -35.765 78.045 -35.720 ;
        RECT 83.165 -35.765 83.545 -35.720 ;
        RECT 77.615 -36.080 83.550 -35.765 ;
        RECT 77.665 -36.100 78.045 -36.080 ;
        RECT 83.165 -36.100 83.545 -36.080 ;
        RECT 87.165 -36.100 87.545 -35.720 ;
        RECT 91.165 -36.100 91.545 -35.720 ;
        RECT 96.875 -35.800 98.615 -35.510 ;
        RECT 100.665 -35.850 101.865 -35.560 ;
        RECT 103.375 -35.890 106.005 -35.435 ;
        RECT 107.585 -35.785 107.965 -35.405 ;
        RECT 61.755 -36.725 82.530 -36.350 ;
        RECT 32.455 -37.225 59.765 -36.885 ;
        RECT 12.070 -37.930 19.330 -37.630 ;
        RECT 12.625 -38.465 16.710 -38.195 ;
        RECT 23.030 -38.230 26.780 -37.955 ;
        RECT 60.785 -38.080 92.750 -37.690 ;
        RECT 105.560 -38.320 108.690 -38.045 ;
        RECT 109.435 -38.080 109.815 -30.920 ;
        RECT 110.675 -33.380 117.415 -33.080 ;
        RECT 111.265 -35.175 114.720 -34.735 ;
        RECT 117.725 -35.335 118.105 -34.955 ;
        RECT 116.125 -35.850 117.325 -35.560 ;
        RECT 123.045 -35.785 123.425 -35.405 ;
        RECT 110.080 -36.560 126.000 -36.260 ;
        RECT 110.615 -37.305 127.560 -37.005 ;
        RECT 28.085 -38.355 46.755 -38.345 ;
        RECT 28.085 -38.435 58.105 -38.355 ;
        RECT 28.085 -38.445 85.190 -38.435 ;
        RECT 28.085 -38.665 94.195 -38.445 ;
        RECT 57.630 -38.755 94.195 -38.665 ;
        RECT -4.015 -44.955 -3.635 -39.125 ;
        RECT 0.240 -40.305 10.895 -39.970 ;
        RECT 0.210 -41.625 1.990 -41.335 ;
        RECT 7.585 -41.655 8.895 -41.335 ;
        RECT -1.060 -42.240 -0.680 -41.860 ;
        RECT 5.395 -42.210 5.775 -41.830 ;
        RECT -3.265 -44.955 0.830 -44.950 ;
        RECT 11.445 -44.955 11.825 -39.125 ;
        RECT 111.810 -39.215 115.940 -38.915 ;
        RECT 27.555 -39.425 63.465 -39.335 ;
        RECT 16.285 -39.725 22.675 -39.435 ;
        RECT 27.555 -39.605 94.595 -39.425 ;
        RECT 62.850 -39.695 94.595 -39.605 ;
        RECT 98.815 -39.815 105.205 -39.525 ;
        RECT 15.700 -40.305 26.205 -39.970 ;
        RECT 51.175 -40.170 61.725 -39.835 ;
        RECT 98.230 -40.395 108.710 -40.060 ;
        RECT 31.770 -40.810 35.070 -40.430 ;
        RECT 35.770 -40.810 39.070 -40.430 ;
        RECT 45.270 -40.810 48.570 -40.430 ;
        RECT 49.270 -40.810 52.570 -40.430 ;
        RECT 68.200 -40.900 69.505 -40.520 ;
        RECT 74.205 -40.900 77.505 -40.520 ;
        RECT 78.205 -40.900 79.565 -40.520 ;
        RECT 81.540 -40.900 83.005 -40.520 ;
        RECT 83.705 -40.900 87.005 -40.520 ;
        RECT 91.705 -40.900 92.885 -40.520 ;
        RECT 31.230 -41.155 31.610 -41.120 ;
        RECT 13.265 -41.640 13.645 -41.260 ;
        RECT 15.670 -41.625 17.450 -41.335 ;
        RECT 18.925 -41.535 20.115 -41.250 ;
        RECT 23.045 -41.655 24.355 -41.335 ;
        RECT 30.965 -41.465 33.975 -41.155 ;
        RECT 31.230 -41.500 31.610 -41.465 ;
        RECT 35.230 -41.500 36.320 -41.120 ;
        RECT 39.230 -41.125 39.610 -41.120 ;
        RECT 36.750 -41.490 39.615 -41.125 ;
        RECT 44.730 -41.145 45.110 -41.120 ;
        RECT 44.715 -41.465 46.860 -41.145 ;
        RECT 39.230 -41.500 39.610 -41.490 ;
        RECT 44.730 -41.500 45.110 -41.465 ;
        RECT 47.775 -41.500 49.110 -41.120 ;
        RECT 52.730 -41.140 53.110 -41.120 ;
        RECT 50.265 -41.460 53.175 -41.140 ;
        RECT 69.665 -41.245 70.045 -41.210 ;
        RECT 52.730 -41.500 53.110 -41.460 ;
        RECT 69.400 -41.555 72.410 -41.245 ;
        RECT 69.665 -41.590 70.045 -41.555 ;
        RECT 73.665 -41.590 74.755 -41.210 ;
        RECT 77.665 -41.215 78.045 -41.210 ;
        RECT 75.185 -41.580 78.050 -41.215 ;
        RECT 83.165 -41.235 83.545 -41.210 ;
        RECT 83.150 -41.555 85.295 -41.235 ;
        RECT 77.665 -41.590 78.045 -41.580 ;
        RECT 83.165 -41.590 83.545 -41.555 ;
        RECT 86.210 -41.590 87.545 -41.210 ;
        RECT 91.165 -41.230 91.545 -41.210 ;
        RECT 88.700 -41.550 91.610 -41.230 ;
        RECT 91.165 -41.590 91.545 -41.550 ;
        RECT 95.795 -41.730 96.175 -41.350 ;
        RECT 98.200 -41.715 99.980 -41.425 ;
        RECT 101.455 -41.625 102.645 -41.340 ;
        RECT 105.575 -41.745 106.885 -41.425 ;
        RECT 14.400 -42.240 14.780 -41.860 ;
        RECT 18.145 -42.200 18.525 -41.820 ;
        RECT 20.855 -42.210 21.235 -41.830 ;
        RECT 22.265 -42.365 25.445 -42.045 ;
        RECT 96.930 -42.330 97.310 -41.950 ;
        RECT 100.675 -42.290 101.055 -41.910 ;
        RECT 103.385 -42.300 103.765 -41.920 ;
        RECT 31.770 -42.810 33.055 -42.430 ;
        RECT 51.085 -42.810 52.570 -42.430 ;
        RECT 104.795 -42.455 107.975 -42.135 ;
        RECT 68.015 -42.900 69.505 -42.520 ;
        RECT 91.705 -42.900 92.780 -42.520 ;
        RECT 31.230 -43.500 32.320 -43.120 ;
        RECT 33.275 -43.490 34.795 -43.130 ;
        RECT 35.715 -43.495 48.565 -43.160 ;
        RECT 52.730 -43.165 53.110 -43.120 ;
        RECT 51.995 -43.465 53.305 -43.165 ;
        RECT 52.730 -43.500 53.110 -43.465 ;
        RECT 69.665 -43.590 70.755 -43.210 ;
        RECT 71.710 -43.580 73.230 -43.220 ;
        RECT 74.150 -43.585 87.000 -43.250 ;
        RECT 91.165 -43.255 91.545 -43.210 ;
        RECT 90.430 -43.555 91.740 -43.255 ;
        RECT 91.165 -43.590 91.545 -43.555 ;
        RECT 28.085 -44.085 61.165 -44.010 ;
        RECT 28.085 -44.360 93.175 -44.085 ;
        RECT 60.225 -44.450 93.175 -44.360 ;
        RECT 94.970 -44.460 99.230 -44.105 ;
        RECT 12.195 -44.955 16.290 -44.950 ;
        RECT -4.385 -44.960 0.830 -44.955 ;
        RECT 11.075 -44.960 16.290 -44.955 ;
        RECT 26.535 -44.960 66.785 -44.955 ;
        RECT -4.385 -45.045 66.785 -44.960 ;
        RECT 93.175 -45.045 98.820 -45.040 ;
        RECT 109.435 -45.045 109.815 -39.215 ;
        RECT 118.315 -39.265 122.815 -38.955 ;
        RECT 114.275 -39.815 120.665 -39.525 ;
        RECT 113.040 -40.980 115.960 -40.680 ;
        RECT 119.505 -40.995 122.875 -40.695 ;
        RECT 111.255 -41.730 111.635 -41.350 ;
        RECT 116.915 -41.625 118.105 -41.340 ;
        RECT 116.135 -42.290 116.515 -41.910 ;
        RECT 120.255 -42.455 123.435 -42.135 ;
        RECT 110.535 -43.540 114.685 -43.270 ;
        RECT 110.185 -45.045 114.280 -45.040 ;
        RECT -4.385 -45.050 98.820 -45.045 ;
        RECT 109.065 -45.050 114.280 -45.045 ;
        RECT -4.385 -45.855 124.095 -45.050 ;
        RECT 66.520 -45.945 124.095 -45.855 ;
        RECT -4.195 -49.665 68.195 -49.640 ;
        RECT -4.195 -50.540 124.250 -49.665 ;
        RECT -3.825 -57.700 -3.445 -50.540 ;
        RECT 1.750 -54.995 2.130 -54.615 ;
        RECT 8.650 -55.005 9.030 -54.625 ;
        RECT -0.925 -55.420 0.815 -55.130 ;
        RECT 5.575 -55.500 8.185 -55.075 ;
        RECT 7.760 -57.940 10.865 -57.665 ;
        RECT 11.635 -57.700 12.015 -50.540 ;
        RECT 67.895 -50.565 124.250 -50.540 ;
        RECT 28.275 -51.550 65.825 -51.525 ;
        RECT 28.275 -51.810 93.655 -51.550 ;
        RECT 64.880 -51.835 93.655 -51.810 ;
        RECT 95.325 -51.855 102.030 -51.555 ;
        RECT 31.980 -52.720 33.180 -52.340 ;
        RECT 34.935 -52.935 37.210 -52.425 ;
        RECT 39.835 -52.935 42.135 -52.425 ;
        RECT 44.430 -52.935 46.710 -52.425 ;
        RECT 51.505 -52.620 52.740 -52.240 ;
        RECT 68.185 -52.745 69.640 -52.365 ;
        RECT 52.920 -52.975 53.300 -52.940 ;
        RECT 73.335 -52.960 75.610 -52.450 ;
        RECT 78.235 -52.960 80.535 -52.450 ;
        RECT 82.830 -52.960 85.110 -52.450 ;
        RECT 91.880 -52.645 93.160 -52.265 ;
        RECT 31.420 -53.080 31.800 -53.040 ;
        RECT 31.350 -53.385 34.185 -53.080 ;
        RECT 50.165 -53.285 53.300 -52.975 ;
        RECT 91.320 -53.000 91.700 -52.965 ;
        RECT 69.820 -53.105 70.200 -53.065 ;
        RECT 52.920 -53.320 53.300 -53.285 ;
        RECT 31.420 -53.420 31.800 -53.385 ;
        RECT 69.750 -53.410 72.585 -53.105 ;
        RECT 88.565 -53.310 91.700 -53.000 ;
        RECT 91.320 -53.345 91.700 -53.310 ;
        RECT 69.820 -53.445 70.200 -53.410 ;
        RECT 13.465 -54.795 16.870 -54.355 ;
        RECT 17.210 -54.995 17.590 -54.615 ;
        RECT 19.925 -54.955 20.305 -54.575 ;
        RECT 24.110 -55.005 24.490 -54.625 ;
        RECT 31.980 -55.020 35.240 -54.640 ;
        RECT 35.980 -55.020 39.240 -54.640 ;
        RECT 45.480 -55.020 48.740 -54.640 ;
        RECT 49.480 -55.020 52.740 -54.640 ;
        RECT 14.535 -55.420 16.275 -55.130 ;
        RECT 18.325 -55.470 19.525 -55.180 ;
        RECT 21.035 -55.500 23.630 -55.125 ;
        RECT 25.245 -55.405 25.625 -55.025 ;
        RECT 68.345 -55.045 69.640 -54.665 ;
        RECT 74.380 -55.045 77.640 -54.665 ;
        RECT 78.380 -55.045 79.565 -54.665 ;
        RECT 81.830 -55.045 83.140 -54.665 ;
        RECT 83.880 -55.045 87.140 -54.665 ;
        RECT 91.880 -55.045 92.895 -54.665 ;
        RECT 95.960 -54.800 99.375 -54.380 ;
        RECT 99.705 -55.020 100.085 -54.640 ;
        RECT 102.420 -54.980 102.800 -54.600 ;
        RECT 106.605 -55.030 106.985 -54.650 ;
        RECT 31.420 -55.720 31.800 -55.340 ;
        RECT 35.420 -55.720 35.800 -55.340 ;
        RECT 39.420 -55.385 39.800 -55.340 ;
        RECT 44.920 -55.385 45.300 -55.340 ;
        RECT 39.370 -55.700 45.305 -55.385 ;
        RECT 39.420 -55.720 39.800 -55.700 ;
        RECT 44.920 -55.720 45.300 -55.700 ;
        RECT 48.920 -55.720 49.300 -55.340 ;
        RECT 52.920 -55.720 53.300 -55.340 ;
        RECT 69.820 -55.745 70.200 -55.365 ;
        RECT 73.820 -55.745 74.200 -55.365 ;
        RECT 77.820 -55.410 78.200 -55.365 ;
        RECT 83.320 -55.410 83.700 -55.365 ;
        RECT 77.770 -55.725 83.705 -55.410 ;
        RECT 77.820 -55.745 78.200 -55.725 ;
        RECT 83.320 -55.745 83.700 -55.725 ;
        RECT 87.320 -55.745 87.700 -55.365 ;
        RECT 91.320 -55.745 91.700 -55.365 ;
        RECT 97.030 -55.445 98.770 -55.155 ;
        RECT 100.820 -55.495 102.020 -55.205 ;
        RECT 103.530 -55.535 106.160 -55.080 ;
        RECT 107.740 -55.430 108.120 -55.050 ;
        RECT 61.910 -56.370 82.685 -55.995 ;
        RECT 32.645 -56.935 59.955 -56.595 ;
        RECT 12.260 -57.640 19.520 -57.340 ;
        RECT 12.815 -58.175 16.900 -57.905 ;
        RECT 23.220 -57.940 26.970 -57.665 ;
        RECT 60.940 -57.725 92.905 -57.335 ;
        RECT 105.715 -57.965 108.845 -57.690 ;
        RECT 109.590 -57.725 109.970 -50.565 ;
        RECT 110.830 -53.025 117.570 -52.725 ;
        RECT 111.420 -54.820 114.875 -54.380 ;
        RECT 117.880 -54.980 118.260 -54.600 ;
        RECT 116.280 -55.495 117.480 -55.205 ;
        RECT 123.200 -55.430 123.580 -55.050 ;
        RECT 110.235 -56.205 126.155 -55.905 ;
        RECT 110.770 -56.950 127.715 -56.650 ;
        RECT 28.275 -58.065 46.945 -58.055 ;
        RECT 28.275 -58.080 58.295 -58.065 ;
        RECT 28.275 -58.090 85.345 -58.080 ;
        RECT 28.275 -58.375 94.350 -58.090 ;
        RECT 57.785 -58.400 94.350 -58.375 ;
        RECT -3.825 -64.665 -3.445 -58.835 ;
        RECT 0.430 -60.015 11.085 -59.680 ;
        RECT 0.400 -61.335 2.180 -61.045 ;
        RECT 7.775 -61.365 9.085 -61.045 ;
        RECT -0.870 -61.950 -0.490 -61.570 ;
        RECT 5.585 -61.920 5.965 -61.540 ;
        RECT -3.075 -64.665 1.020 -64.660 ;
        RECT 11.635 -64.665 12.015 -58.835 ;
        RECT 111.965 -58.860 116.095 -58.560 ;
        RECT 27.745 -59.070 63.655 -59.045 ;
        RECT 16.475 -59.435 22.865 -59.145 ;
        RECT 27.745 -59.315 94.750 -59.070 ;
        RECT 63.005 -59.340 94.750 -59.315 ;
        RECT 98.970 -59.460 105.360 -59.170 ;
        RECT 15.890 -60.015 26.395 -59.680 ;
        RECT 51.365 -59.880 61.915 -59.545 ;
        RECT 98.385 -60.040 108.865 -59.705 ;
        RECT 31.960 -60.520 35.260 -60.140 ;
        RECT 35.960 -60.520 39.260 -60.140 ;
        RECT 45.460 -60.520 48.760 -60.140 ;
        RECT 49.460 -60.520 52.760 -60.140 ;
        RECT 68.355 -60.545 69.660 -60.165 ;
        RECT 74.360 -60.545 77.660 -60.165 ;
        RECT 78.360 -60.545 79.720 -60.165 ;
        RECT 81.695 -60.545 83.160 -60.165 ;
        RECT 83.860 -60.545 87.160 -60.165 ;
        RECT 91.860 -60.545 93.040 -60.165 ;
        RECT 31.420 -60.865 31.800 -60.830 ;
        RECT 13.455 -61.350 13.835 -60.970 ;
        RECT 15.860 -61.335 17.640 -61.045 ;
        RECT 19.115 -61.245 20.305 -60.960 ;
        RECT 23.235 -61.365 24.545 -61.045 ;
        RECT 31.155 -61.175 34.165 -60.865 ;
        RECT 31.420 -61.210 31.800 -61.175 ;
        RECT 35.420 -61.210 36.510 -60.830 ;
        RECT 39.420 -60.835 39.800 -60.830 ;
        RECT 36.940 -61.200 39.805 -60.835 ;
        RECT 44.920 -60.855 45.300 -60.830 ;
        RECT 44.905 -61.175 47.050 -60.855 ;
        RECT 39.420 -61.210 39.800 -61.200 ;
        RECT 44.920 -61.210 45.300 -61.175 ;
        RECT 47.965 -61.210 49.300 -60.830 ;
        RECT 52.920 -60.850 53.300 -60.830 ;
        RECT 50.455 -61.170 53.365 -60.850 ;
        RECT 69.820 -60.890 70.200 -60.855 ;
        RECT 52.920 -61.210 53.300 -61.170 ;
        RECT 69.555 -61.200 72.565 -60.890 ;
        RECT 69.820 -61.235 70.200 -61.200 ;
        RECT 73.820 -61.235 74.910 -60.855 ;
        RECT 77.820 -60.860 78.200 -60.855 ;
        RECT 75.340 -61.225 78.205 -60.860 ;
        RECT 83.320 -60.880 83.700 -60.855 ;
        RECT 83.305 -61.200 85.450 -60.880 ;
        RECT 77.820 -61.235 78.200 -61.225 ;
        RECT 83.320 -61.235 83.700 -61.200 ;
        RECT 86.365 -61.235 87.700 -60.855 ;
        RECT 91.320 -60.875 91.700 -60.855 ;
        RECT 88.855 -61.195 91.765 -60.875 ;
        RECT 91.320 -61.235 91.700 -61.195 ;
        RECT 95.950 -61.375 96.330 -60.995 ;
        RECT 98.355 -61.360 100.135 -61.070 ;
        RECT 101.610 -61.270 102.800 -60.985 ;
        RECT 105.730 -61.390 107.040 -61.070 ;
        RECT 14.590 -61.950 14.970 -61.570 ;
        RECT 18.335 -61.910 18.715 -61.530 ;
        RECT 21.045 -61.920 21.425 -61.540 ;
        RECT 22.455 -62.075 25.635 -61.755 ;
        RECT 97.085 -61.975 97.465 -61.595 ;
        RECT 100.830 -61.935 101.210 -61.555 ;
        RECT 103.540 -61.945 103.920 -61.565 ;
        RECT 104.950 -62.100 108.130 -61.780 ;
        RECT 31.960 -62.520 33.245 -62.140 ;
        RECT 51.275 -62.520 52.760 -62.140 ;
        RECT 68.170 -62.545 69.660 -62.165 ;
        RECT 91.860 -62.545 92.935 -62.165 ;
        RECT 31.420 -63.210 32.510 -62.830 ;
        RECT 33.465 -63.200 34.985 -62.840 ;
        RECT 35.905 -63.205 48.755 -62.870 ;
        RECT 52.920 -62.875 53.300 -62.830 ;
        RECT 52.185 -63.175 53.495 -62.875 ;
        RECT 52.920 -63.210 53.300 -63.175 ;
        RECT 69.820 -63.235 70.910 -62.855 ;
        RECT 71.865 -63.225 73.385 -62.865 ;
        RECT 74.305 -63.230 87.155 -62.895 ;
        RECT 91.320 -62.900 91.700 -62.855 ;
        RECT 90.585 -63.200 91.895 -62.900 ;
        RECT 91.320 -63.235 91.700 -63.200 ;
        RECT 28.275 -63.730 61.355 -63.720 ;
        RECT 28.275 -64.070 93.330 -63.730 ;
        RECT 60.380 -64.095 93.330 -64.070 ;
        RECT 95.125 -64.105 99.385 -63.750 ;
        RECT 12.385 -64.665 16.480 -64.660 ;
        RECT -4.195 -64.670 1.020 -64.665 ;
        RECT 11.265 -64.670 16.480 -64.665 ;
        RECT 26.725 -64.670 66.975 -64.665 ;
        RECT -4.195 -64.690 66.975 -64.670 ;
        RECT 93.330 -64.690 98.975 -64.685 ;
        RECT 109.590 -64.690 109.970 -58.860 ;
        RECT 118.470 -58.910 122.970 -58.600 ;
        RECT 114.430 -59.460 120.820 -59.170 ;
        RECT 113.195 -60.625 116.115 -60.325 ;
        RECT 119.660 -60.640 123.030 -60.340 ;
        RECT 111.410 -61.375 111.790 -60.995 ;
        RECT 117.070 -61.270 118.260 -60.985 ;
        RECT 116.290 -61.935 116.670 -61.555 ;
        RECT 120.410 -62.100 123.590 -61.780 ;
        RECT 110.690 -63.185 114.840 -62.915 ;
        RECT 110.340 -64.690 114.435 -64.685 ;
        RECT -4.195 -64.695 98.975 -64.690 ;
        RECT 109.220 -64.695 114.435 -64.690 ;
        RECT -4.195 -65.565 124.250 -64.695 ;
        RECT 66.675 -65.590 124.250 -65.565 ;
        RECT 67.895 -69.480 124.250 -69.460 ;
        RECT -4.390 -70.360 124.250 -69.480 ;
        RECT -4.390 -70.380 68.000 -70.360 ;
        RECT -4.020 -77.540 -3.640 -70.380 ;
        RECT 1.555 -74.835 1.935 -74.455 ;
        RECT 8.455 -74.845 8.835 -74.465 ;
        RECT -1.120 -75.260 0.620 -74.970 ;
        RECT 5.380 -75.340 7.990 -74.915 ;
        RECT 7.565 -77.780 10.670 -77.505 ;
        RECT 11.440 -77.540 11.820 -70.380 ;
        RECT 64.880 -71.365 93.655 -71.345 ;
        RECT 28.080 -71.630 93.655 -71.365 ;
        RECT 28.080 -71.650 65.630 -71.630 ;
        RECT 95.325 -71.650 102.030 -71.350 ;
        RECT 31.785 -72.560 32.985 -72.180 ;
        RECT 34.740 -72.775 37.015 -72.265 ;
        RECT 39.640 -72.775 41.940 -72.265 ;
        RECT 44.235 -72.775 46.515 -72.265 ;
        RECT 51.310 -72.460 52.545 -72.080 ;
        RECT 68.185 -72.540 69.640 -72.160 ;
        RECT 73.335 -72.755 75.610 -72.245 ;
        RECT 78.235 -72.755 80.535 -72.245 ;
        RECT 82.830 -72.755 85.110 -72.245 ;
        RECT 91.880 -72.440 93.160 -72.060 ;
        RECT 52.725 -72.815 53.105 -72.780 ;
        RECT 91.320 -72.795 91.700 -72.760 ;
        RECT 31.225 -72.920 31.605 -72.880 ;
        RECT 31.155 -73.225 33.990 -72.920 ;
        RECT 49.970 -73.125 53.105 -72.815 ;
        RECT 69.820 -72.900 70.200 -72.860 ;
        RECT 52.725 -73.160 53.105 -73.125 ;
        RECT 69.750 -73.205 72.585 -72.900 ;
        RECT 88.565 -73.105 91.700 -72.795 ;
        RECT 91.320 -73.140 91.700 -73.105 ;
        RECT 31.225 -73.260 31.605 -73.225 ;
        RECT 69.820 -73.240 70.200 -73.205 ;
        RECT 13.270 -74.635 16.675 -74.195 ;
        RECT 17.015 -74.835 17.395 -74.455 ;
        RECT 19.730 -74.795 20.110 -74.415 ;
        RECT 23.915 -74.845 24.295 -74.465 ;
        RECT 31.785 -74.860 35.045 -74.480 ;
        RECT 35.785 -74.860 39.045 -74.480 ;
        RECT 45.285 -74.860 48.545 -74.480 ;
        RECT 49.285 -74.860 52.545 -74.480 ;
        RECT 68.345 -74.840 69.640 -74.460 ;
        RECT 74.380 -74.840 77.640 -74.460 ;
        RECT 78.380 -74.840 79.565 -74.460 ;
        RECT 81.830 -74.840 83.140 -74.460 ;
        RECT 83.880 -74.840 87.140 -74.460 ;
        RECT 91.880 -74.840 92.895 -74.460 ;
        RECT 95.960 -74.595 99.375 -74.175 ;
        RECT 99.705 -74.815 100.085 -74.435 ;
        RECT 102.420 -74.775 102.800 -74.395 ;
        RECT 106.605 -74.825 106.985 -74.445 ;
        RECT 14.340 -75.260 16.080 -74.970 ;
        RECT 18.130 -75.310 19.330 -75.020 ;
        RECT 20.840 -75.340 23.435 -74.965 ;
        RECT 25.050 -75.245 25.430 -74.865 ;
        RECT 31.225 -75.560 31.605 -75.180 ;
        RECT 35.225 -75.560 35.605 -75.180 ;
        RECT 39.225 -75.225 39.605 -75.180 ;
        RECT 44.725 -75.225 45.105 -75.180 ;
        RECT 39.175 -75.540 45.110 -75.225 ;
        RECT 39.225 -75.560 39.605 -75.540 ;
        RECT 44.725 -75.560 45.105 -75.540 ;
        RECT 48.725 -75.560 49.105 -75.180 ;
        RECT 52.725 -75.560 53.105 -75.180 ;
        RECT 69.820 -75.540 70.200 -75.160 ;
        RECT 73.820 -75.540 74.200 -75.160 ;
        RECT 77.820 -75.205 78.200 -75.160 ;
        RECT 83.320 -75.205 83.700 -75.160 ;
        RECT 77.770 -75.520 83.705 -75.205 ;
        RECT 77.820 -75.540 78.200 -75.520 ;
        RECT 83.320 -75.540 83.700 -75.520 ;
        RECT 87.320 -75.540 87.700 -75.160 ;
        RECT 91.320 -75.540 91.700 -75.160 ;
        RECT 97.030 -75.240 98.770 -74.950 ;
        RECT 100.820 -75.290 102.020 -75.000 ;
        RECT 103.530 -75.330 106.160 -74.875 ;
        RECT 107.740 -75.225 108.120 -74.845 ;
        RECT 61.910 -76.165 82.685 -75.790 ;
        RECT 32.450 -76.775 59.760 -76.435 ;
        RECT 12.065 -77.480 19.325 -77.180 ;
        RECT 12.620 -78.015 16.705 -77.745 ;
        RECT 23.025 -77.780 26.775 -77.505 ;
        RECT 60.940 -77.520 92.905 -77.130 ;
        RECT 105.715 -77.760 108.845 -77.485 ;
        RECT 109.590 -77.520 109.970 -70.360 ;
        RECT 110.830 -72.820 117.570 -72.520 ;
        RECT 111.420 -74.615 114.875 -74.175 ;
        RECT 117.880 -74.775 118.260 -74.395 ;
        RECT 116.280 -75.290 117.480 -75.000 ;
        RECT 123.200 -75.225 123.580 -74.845 ;
        RECT 110.235 -76.000 126.155 -75.700 ;
        RECT 110.770 -76.745 127.715 -76.445 ;
        RECT 57.785 -77.885 85.345 -77.875 ;
        RECT 28.080 -77.905 46.750 -77.895 ;
        RECT 57.785 -77.905 94.350 -77.885 ;
        RECT 28.080 -78.195 94.350 -77.905 ;
        RECT 28.080 -78.215 58.100 -78.195 ;
        RECT 111.965 -78.655 116.095 -78.355 ;
        RECT -4.020 -84.505 -3.640 -78.675 ;
        RECT 0.235 -79.855 10.890 -79.520 ;
        RECT 0.205 -81.175 1.985 -80.885 ;
        RECT 7.580 -81.205 8.890 -80.885 ;
        RECT -1.065 -81.790 -0.685 -81.410 ;
        RECT 5.390 -81.760 5.770 -81.380 ;
        RECT -3.270 -84.505 0.825 -84.500 ;
        RECT 11.440 -84.505 11.820 -78.675 ;
        RECT 63.005 -78.885 94.750 -78.865 ;
        RECT 16.280 -79.275 22.670 -78.985 ;
        RECT 27.550 -79.135 94.750 -78.885 ;
        RECT 27.550 -79.155 63.460 -79.135 ;
        RECT 98.970 -79.255 105.360 -78.965 ;
        RECT 15.695 -79.855 26.200 -79.520 ;
        RECT 51.170 -79.720 61.720 -79.385 ;
        RECT 98.385 -79.835 108.865 -79.500 ;
        RECT 31.765 -80.360 35.065 -79.980 ;
        RECT 35.765 -80.360 39.065 -79.980 ;
        RECT 45.265 -80.360 48.565 -79.980 ;
        RECT 49.265 -80.360 52.565 -79.980 ;
        RECT 68.355 -80.340 69.660 -79.960 ;
        RECT 74.360 -80.340 77.660 -79.960 ;
        RECT 78.360 -80.340 79.720 -79.960 ;
        RECT 81.695 -80.340 83.160 -79.960 ;
        RECT 83.860 -80.340 87.160 -79.960 ;
        RECT 91.860 -80.340 93.040 -79.960 ;
        RECT 31.225 -80.705 31.605 -80.670 ;
        RECT 13.260 -81.190 13.640 -80.810 ;
        RECT 15.665 -81.175 17.445 -80.885 ;
        RECT 18.920 -81.085 20.110 -80.800 ;
        RECT 23.040 -81.205 24.350 -80.885 ;
        RECT 30.960 -81.015 33.970 -80.705 ;
        RECT 31.225 -81.050 31.605 -81.015 ;
        RECT 35.225 -81.050 36.315 -80.670 ;
        RECT 39.225 -80.675 39.605 -80.670 ;
        RECT 36.745 -81.040 39.610 -80.675 ;
        RECT 44.725 -80.695 45.105 -80.670 ;
        RECT 44.710 -81.015 46.855 -80.695 ;
        RECT 39.225 -81.050 39.605 -81.040 ;
        RECT 44.725 -81.050 45.105 -81.015 ;
        RECT 47.770 -81.050 49.105 -80.670 ;
        RECT 52.725 -80.690 53.105 -80.670 ;
        RECT 69.820 -80.685 70.200 -80.650 ;
        RECT 50.260 -81.010 53.170 -80.690 ;
        RECT 69.555 -80.995 72.565 -80.685 ;
        RECT 52.725 -81.050 53.105 -81.010 ;
        RECT 69.820 -81.030 70.200 -80.995 ;
        RECT 73.820 -81.030 74.910 -80.650 ;
        RECT 77.820 -80.655 78.200 -80.650 ;
        RECT 75.340 -81.020 78.205 -80.655 ;
        RECT 83.320 -80.675 83.700 -80.650 ;
        RECT 83.305 -80.995 85.450 -80.675 ;
        RECT 77.820 -81.030 78.200 -81.020 ;
        RECT 83.320 -81.030 83.700 -80.995 ;
        RECT 86.365 -81.030 87.700 -80.650 ;
        RECT 91.320 -80.670 91.700 -80.650 ;
        RECT 88.855 -80.990 91.765 -80.670 ;
        RECT 91.320 -81.030 91.700 -80.990 ;
        RECT 95.950 -81.170 96.330 -80.790 ;
        RECT 98.355 -81.155 100.135 -80.865 ;
        RECT 101.610 -81.065 102.800 -80.780 ;
        RECT 105.730 -81.185 107.040 -80.865 ;
        RECT 14.395 -81.790 14.775 -81.410 ;
        RECT 18.140 -81.750 18.520 -81.370 ;
        RECT 20.850 -81.760 21.230 -81.380 ;
        RECT 22.260 -81.915 25.440 -81.595 ;
        RECT 97.085 -81.770 97.465 -81.390 ;
        RECT 100.830 -81.730 101.210 -81.350 ;
        RECT 103.540 -81.740 103.920 -81.360 ;
        RECT 104.950 -81.895 108.130 -81.575 ;
        RECT 31.765 -82.360 33.050 -81.980 ;
        RECT 51.080 -82.360 52.565 -81.980 ;
        RECT 68.170 -82.340 69.660 -81.960 ;
        RECT 91.860 -82.340 92.935 -81.960 ;
        RECT 31.225 -83.050 32.315 -82.670 ;
        RECT 33.270 -83.040 34.790 -82.680 ;
        RECT 35.710 -83.045 48.560 -82.710 ;
        RECT 52.725 -82.715 53.105 -82.670 ;
        RECT 51.990 -83.015 53.300 -82.715 ;
        RECT 52.725 -83.050 53.105 -83.015 ;
        RECT 69.820 -83.030 70.910 -82.650 ;
        RECT 71.865 -83.020 73.385 -82.660 ;
        RECT 74.305 -83.025 87.155 -82.690 ;
        RECT 91.320 -82.695 91.700 -82.650 ;
        RECT 90.585 -82.995 91.895 -82.695 ;
        RECT 91.320 -83.030 91.700 -82.995 ;
        RECT 60.380 -83.560 93.330 -83.525 ;
        RECT 28.080 -83.890 93.330 -83.560 ;
        RECT 28.080 -83.910 61.160 -83.890 ;
        RECT 95.125 -83.900 99.385 -83.545 ;
        RECT 93.330 -84.485 98.975 -84.480 ;
        RECT 109.590 -84.485 109.970 -78.655 ;
        RECT 118.470 -78.705 122.970 -78.395 ;
        RECT 114.430 -79.255 120.820 -78.965 ;
        RECT 113.195 -80.420 116.115 -80.120 ;
        RECT 119.660 -80.435 123.030 -80.135 ;
        RECT 111.410 -81.170 111.790 -80.790 ;
        RECT 117.070 -81.065 118.260 -80.780 ;
        RECT 116.290 -81.730 116.670 -81.350 ;
        RECT 120.410 -81.895 123.590 -81.575 ;
        RECT 110.690 -82.980 114.840 -82.710 ;
        RECT 110.340 -84.485 114.435 -84.480 ;
        RECT 66.675 -84.490 98.975 -84.485 ;
        RECT 109.220 -84.490 114.435 -84.485 ;
        RECT 12.190 -84.505 16.285 -84.500 ;
        RECT 66.675 -84.505 124.250 -84.490 ;
        RECT -4.390 -84.510 0.825 -84.505 ;
        RECT 11.070 -84.510 16.285 -84.505 ;
        RECT 26.530 -84.510 124.250 -84.505 ;
        RECT -4.390 -85.385 124.250 -84.510 ;
        RECT -4.390 -85.405 66.780 -85.385 ;
        RECT -4.520 -89.215 67.870 -89.190 ;
        RECT -4.520 -90.090 124.170 -89.215 ;
        RECT -4.150 -97.250 -3.770 -90.090 ;
        RECT 1.425 -94.545 1.805 -94.165 ;
        RECT 8.325 -94.555 8.705 -94.175 ;
        RECT -1.250 -94.970 0.490 -94.680 ;
        RECT 5.250 -95.050 7.860 -94.625 ;
        RECT 7.435 -97.490 10.540 -97.215 ;
        RECT 11.310 -97.250 11.690 -90.090 ;
        RECT 67.815 -90.115 124.170 -90.090 ;
        RECT 27.950 -91.100 65.500 -91.075 ;
        RECT 27.950 -91.360 93.575 -91.100 ;
        RECT 64.800 -91.385 93.575 -91.360 ;
        RECT 95.245 -91.405 101.950 -91.105 ;
        RECT 31.655 -92.270 32.855 -91.890 ;
        RECT 34.610 -92.485 36.885 -91.975 ;
        RECT 39.510 -92.485 41.810 -91.975 ;
        RECT 44.105 -92.485 46.385 -91.975 ;
        RECT 51.180 -92.170 52.415 -91.790 ;
        RECT 68.105 -92.295 69.560 -91.915 ;
        RECT 52.595 -92.525 52.975 -92.490 ;
        RECT 73.255 -92.510 75.530 -92.000 ;
        RECT 78.155 -92.510 80.455 -92.000 ;
        RECT 82.750 -92.510 85.030 -92.000 ;
        RECT 91.800 -92.195 93.080 -91.815 ;
        RECT 31.095 -92.630 31.475 -92.590 ;
        RECT 31.025 -92.935 33.860 -92.630 ;
        RECT 49.840 -92.835 52.975 -92.525 ;
        RECT 91.240 -92.550 91.620 -92.515 ;
        RECT 69.740 -92.655 70.120 -92.615 ;
        RECT 52.595 -92.870 52.975 -92.835 ;
        RECT 31.095 -92.970 31.475 -92.935 ;
        RECT 69.670 -92.960 72.505 -92.655 ;
        RECT 88.485 -92.860 91.620 -92.550 ;
        RECT 91.240 -92.895 91.620 -92.860 ;
        RECT 69.740 -92.995 70.120 -92.960 ;
        RECT 13.140 -94.345 16.545 -93.905 ;
        RECT 16.885 -94.545 17.265 -94.165 ;
        RECT 19.600 -94.505 19.980 -94.125 ;
        RECT 23.785 -94.555 24.165 -94.175 ;
        RECT 31.655 -94.570 34.915 -94.190 ;
        RECT 35.655 -94.570 38.915 -94.190 ;
        RECT 45.155 -94.570 48.415 -94.190 ;
        RECT 49.155 -94.570 52.415 -94.190 ;
        RECT 14.210 -94.970 15.950 -94.680 ;
        RECT 18.000 -95.020 19.200 -94.730 ;
        RECT 20.710 -95.050 23.305 -94.675 ;
        RECT 24.920 -94.955 25.300 -94.575 ;
        RECT 68.265 -94.595 69.560 -94.215 ;
        RECT 74.300 -94.595 77.560 -94.215 ;
        RECT 78.300 -94.595 79.485 -94.215 ;
        RECT 81.750 -94.595 83.060 -94.215 ;
        RECT 83.800 -94.595 87.060 -94.215 ;
        RECT 91.800 -94.595 92.815 -94.215 ;
        RECT 95.880 -94.350 99.295 -93.930 ;
        RECT 99.625 -94.570 100.005 -94.190 ;
        RECT 102.340 -94.530 102.720 -94.150 ;
        RECT 106.525 -94.580 106.905 -94.200 ;
        RECT 31.095 -95.270 31.475 -94.890 ;
        RECT 35.095 -95.270 35.475 -94.890 ;
        RECT 39.095 -94.935 39.475 -94.890 ;
        RECT 44.595 -94.935 44.975 -94.890 ;
        RECT 39.045 -95.250 44.980 -94.935 ;
        RECT 39.095 -95.270 39.475 -95.250 ;
        RECT 44.595 -95.270 44.975 -95.250 ;
        RECT 48.595 -95.270 48.975 -94.890 ;
        RECT 52.595 -95.270 52.975 -94.890 ;
        RECT 69.740 -95.295 70.120 -94.915 ;
        RECT 73.740 -95.295 74.120 -94.915 ;
        RECT 77.740 -94.960 78.120 -94.915 ;
        RECT 83.240 -94.960 83.620 -94.915 ;
        RECT 77.690 -95.275 83.625 -94.960 ;
        RECT 77.740 -95.295 78.120 -95.275 ;
        RECT 83.240 -95.295 83.620 -95.275 ;
        RECT 87.240 -95.295 87.620 -94.915 ;
        RECT 91.240 -95.295 91.620 -94.915 ;
        RECT 96.950 -94.995 98.690 -94.705 ;
        RECT 100.740 -95.045 101.940 -94.755 ;
        RECT 103.450 -95.085 106.080 -94.630 ;
        RECT 107.660 -94.980 108.040 -94.600 ;
        RECT 61.830 -95.920 82.605 -95.545 ;
        RECT 32.320 -96.485 59.630 -96.145 ;
        RECT 11.935 -97.190 19.195 -96.890 ;
        RECT 12.490 -97.725 16.575 -97.455 ;
        RECT 22.895 -97.490 26.645 -97.215 ;
        RECT 60.860 -97.275 92.825 -96.885 ;
        RECT 105.635 -97.515 108.765 -97.240 ;
        RECT 109.510 -97.275 109.890 -90.115 ;
        RECT 110.750 -92.575 117.490 -92.275 ;
        RECT 111.340 -94.370 114.795 -93.930 ;
        RECT 117.800 -94.530 118.180 -94.150 ;
        RECT 116.200 -95.045 117.400 -94.755 ;
        RECT 123.120 -94.980 123.500 -94.600 ;
        RECT 110.155 -95.755 126.075 -95.455 ;
        RECT 110.690 -96.500 127.635 -96.200 ;
        RECT 27.950 -97.615 46.620 -97.605 ;
        RECT 27.950 -97.630 57.970 -97.615 ;
        RECT 27.950 -97.640 85.265 -97.630 ;
        RECT 27.950 -97.925 94.270 -97.640 ;
        RECT 57.705 -97.950 94.270 -97.925 ;
        RECT -4.150 -104.215 -3.770 -98.385 ;
        RECT 0.105 -99.565 10.760 -99.230 ;
        RECT 0.075 -100.885 1.855 -100.595 ;
        RECT 7.450 -100.915 8.760 -100.595 ;
        RECT -1.195 -101.500 -0.815 -101.120 ;
        RECT 5.260 -101.470 5.640 -101.090 ;
        RECT -3.400 -104.215 0.695 -104.210 ;
        RECT 11.310 -104.215 11.690 -98.385 ;
        RECT 111.885 -98.410 116.015 -98.110 ;
        RECT 27.420 -98.620 63.330 -98.595 ;
        RECT 16.150 -98.985 22.540 -98.695 ;
        RECT 27.420 -98.865 94.670 -98.620 ;
        RECT 62.925 -98.890 94.670 -98.865 ;
        RECT 98.890 -99.010 105.280 -98.720 ;
        RECT 15.565 -99.565 26.070 -99.230 ;
        RECT 51.040 -99.430 61.590 -99.095 ;
        RECT 98.305 -99.590 108.785 -99.255 ;
        RECT 31.635 -100.070 34.935 -99.690 ;
        RECT 35.635 -100.070 38.935 -99.690 ;
        RECT 45.135 -100.070 48.435 -99.690 ;
        RECT 49.135 -100.070 52.435 -99.690 ;
        RECT 68.275 -100.095 69.580 -99.715 ;
        RECT 74.280 -100.095 77.580 -99.715 ;
        RECT 78.280 -100.095 79.640 -99.715 ;
        RECT 81.615 -100.095 83.080 -99.715 ;
        RECT 83.780 -100.095 87.080 -99.715 ;
        RECT 91.780 -100.095 92.960 -99.715 ;
        RECT 31.095 -100.415 31.475 -100.380 ;
        RECT 13.130 -100.900 13.510 -100.520 ;
        RECT 15.535 -100.885 17.315 -100.595 ;
        RECT 18.790 -100.795 19.980 -100.510 ;
        RECT 22.910 -100.915 24.220 -100.595 ;
        RECT 30.830 -100.725 33.840 -100.415 ;
        RECT 31.095 -100.760 31.475 -100.725 ;
        RECT 35.095 -100.760 36.185 -100.380 ;
        RECT 39.095 -100.385 39.475 -100.380 ;
        RECT 36.615 -100.750 39.480 -100.385 ;
        RECT 44.595 -100.405 44.975 -100.380 ;
        RECT 44.580 -100.725 46.725 -100.405 ;
        RECT 39.095 -100.760 39.475 -100.750 ;
        RECT 44.595 -100.760 44.975 -100.725 ;
        RECT 47.640 -100.760 48.975 -100.380 ;
        RECT 52.595 -100.400 52.975 -100.380 ;
        RECT 50.130 -100.720 53.040 -100.400 ;
        RECT 69.740 -100.440 70.120 -100.405 ;
        RECT 52.595 -100.760 52.975 -100.720 ;
        RECT 69.475 -100.750 72.485 -100.440 ;
        RECT 69.740 -100.785 70.120 -100.750 ;
        RECT 73.740 -100.785 74.830 -100.405 ;
        RECT 77.740 -100.410 78.120 -100.405 ;
        RECT 75.260 -100.775 78.125 -100.410 ;
        RECT 83.240 -100.430 83.620 -100.405 ;
        RECT 83.225 -100.750 85.370 -100.430 ;
        RECT 77.740 -100.785 78.120 -100.775 ;
        RECT 83.240 -100.785 83.620 -100.750 ;
        RECT 86.285 -100.785 87.620 -100.405 ;
        RECT 91.240 -100.425 91.620 -100.405 ;
        RECT 88.775 -100.745 91.685 -100.425 ;
        RECT 91.240 -100.785 91.620 -100.745 ;
        RECT 95.870 -100.925 96.250 -100.545 ;
        RECT 98.275 -100.910 100.055 -100.620 ;
        RECT 101.530 -100.820 102.720 -100.535 ;
        RECT 105.650 -100.940 106.960 -100.620 ;
        RECT 14.265 -101.500 14.645 -101.120 ;
        RECT 18.010 -101.460 18.390 -101.080 ;
        RECT 20.720 -101.470 21.100 -101.090 ;
        RECT 22.130 -101.625 25.310 -101.305 ;
        RECT 97.005 -101.525 97.385 -101.145 ;
        RECT 100.750 -101.485 101.130 -101.105 ;
        RECT 103.460 -101.495 103.840 -101.115 ;
        RECT 104.870 -101.650 108.050 -101.330 ;
        RECT 31.635 -102.070 32.920 -101.690 ;
        RECT 50.950 -102.070 52.435 -101.690 ;
        RECT 68.090 -102.095 69.580 -101.715 ;
        RECT 91.780 -102.095 92.855 -101.715 ;
        RECT 31.095 -102.760 32.185 -102.380 ;
        RECT 33.140 -102.750 34.660 -102.390 ;
        RECT 35.580 -102.755 48.430 -102.420 ;
        RECT 52.595 -102.425 52.975 -102.380 ;
        RECT 51.860 -102.725 53.170 -102.425 ;
        RECT 52.595 -102.760 52.975 -102.725 ;
        RECT 69.740 -102.785 70.830 -102.405 ;
        RECT 71.785 -102.775 73.305 -102.415 ;
        RECT 74.225 -102.780 87.075 -102.445 ;
        RECT 91.240 -102.450 91.620 -102.405 ;
        RECT 90.505 -102.750 91.815 -102.450 ;
        RECT 91.240 -102.785 91.620 -102.750 ;
        RECT 27.950 -103.280 61.030 -103.270 ;
        RECT 27.950 -103.620 93.250 -103.280 ;
        RECT 60.300 -103.645 93.250 -103.620 ;
        RECT 95.045 -103.655 99.305 -103.300 ;
        RECT 12.060 -104.215 16.155 -104.210 ;
        RECT -4.520 -104.220 0.695 -104.215 ;
        RECT 10.940 -104.220 16.155 -104.215 ;
        RECT 26.400 -104.220 66.650 -104.215 ;
        RECT -4.520 -104.240 66.650 -104.220 ;
        RECT 93.250 -104.240 98.895 -104.235 ;
        RECT 109.510 -104.240 109.890 -98.410 ;
        RECT 118.390 -98.460 122.890 -98.150 ;
        RECT 114.350 -99.010 120.740 -98.720 ;
        RECT 113.115 -100.175 116.035 -99.875 ;
        RECT 119.580 -100.190 122.950 -99.890 ;
        RECT 111.330 -100.925 111.710 -100.545 ;
        RECT 116.990 -100.820 118.180 -100.535 ;
        RECT 116.210 -101.485 116.590 -101.105 ;
        RECT 120.330 -101.650 123.510 -101.330 ;
        RECT 110.610 -102.735 114.760 -102.465 ;
        RECT 110.260 -104.240 114.355 -104.235 ;
        RECT -4.520 -104.245 98.895 -104.240 ;
        RECT 109.140 -104.245 114.355 -104.240 ;
        RECT -4.520 -105.115 124.170 -104.245 ;
        RECT 66.595 -105.140 124.170 -105.115 ;
        RECT 67.920 -108.950 124.275 -108.930 ;
        RECT -4.390 -109.830 124.275 -108.950 ;
        RECT -4.390 -109.850 68.000 -109.830 ;
        RECT -4.020 -117.010 -3.640 -109.850 ;
        RECT 1.555 -114.305 1.935 -113.925 ;
        RECT 8.455 -114.315 8.835 -113.935 ;
        RECT -1.120 -114.730 0.620 -114.440 ;
        RECT 5.380 -114.810 7.990 -114.385 ;
        RECT 7.565 -117.250 10.670 -116.975 ;
        RECT 11.440 -117.010 11.820 -109.850 ;
        RECT 64.905 -110.835 93.680 -110.815 ;
        RECT 28.080 -111.100 93.680 -110.835 ;
        RECT 28.080 -111.120 65.630 -111.100 ;
        RECT 95.350 -111.120 102.055 -110.820 ;
        RECT 31.785 -112.030 32.985 -111.650 ;
        RECT 34.740 -112.245 37.015 -111.735 ;
        RECT 39.640 -112.245 41.940 -111.735 ;
        RECT 44.235 -112.245 46.515 -111.735 ;
        RECT 51.310 -111.930 52.545 -111.550 ;
        RECT 68.210 -112.010 69.665 -111.630 ;
        RECT 73.360 -112.225 75.635 -111.715 ;
        RECT 78.260 -112.225 80.560 -111.715 ;
        RECT 82.855 -112.225 85.135 -111.715 ;
        RECT 91.905 -111.910 93.185 -111.530 ;
        RECT 52.725 -112.285 53.105 -112.250 ;
        RECT 91.345 -112.265 91.725 -112.230 ;
        RECT 31.225 -112.390 31.605 -112.350 ;
        RECT 31.155 -112.695 33.990 -112.390 ;
        RECT 49.970 -112.595 53.105 -112.285 ;
        RECT 69.845 -112.370 70.225 -112.330 ;
        RECT 52.725 -112.630 53.105 -112.595 ;
        RECT 69.775 -112.675 72.610 -112.370 ;
        RECT 88.590 -112.575 91.725 -112.265 ;
        RECT 91.345 -112.610 91.725 -112.575 ;
        RECT 31.225 -112.730 31.605 -112.695 ;
        RECT 69.845 -112.710 70.225 -112.675 ;
        RECT 13.270 -114.105 16.675 -113.665 ;
        RECT 17.015 -114.305 17.395 -113.925 ;
        RECT 19.730 -114.265 20.110 -113.885 ;
        RECT 23.915 -114.315 24.295 -113.935 ;
        RECT 31.785 -114.330 35.045 -113.950 ;
        RECT 35.785 -114.330 39.045 -113.950 ;
        RECT 45.285 -114.330 48.545 -113.950 ;
        RECT 49.285 -114.330 52.545 -113.950 ;
        RECT 68.370 -114.310 69.665 -113.930 ;
        RECT 74.405 -114.310 77.665 -113.930 ;
        RECT 78.405 -114.310 79.590 -113.930 ;
        RECT 81.855 -114.310 83.165 -113.930 ;
        RECT 83.905 -114.310 87.165 -113.930 ;
        RECT 91.905 -114.310 92.920 -113.930 ;
        RECT 95.985 -114.065 99.400 -113.645 ;
        RECT 99.730 -114.285 100.110 -113.905 ;
        RECT 102.445 -114.245 102.825 -113.865 ;
        RECT 106.630 -114.295 107.010 -113.915 ;
        RECT 14.340 -114.730 16.080 -114.440 ;
        RECT 18.130 -114.780 19.330 -114.490 ;
        RECT 20.840 -114.810 23.435 -114.435 ;
        RECT 25.050 -114.715 25.430 -114.335 ;
        RECT 31.225 -115.030 31.605 -114.650 ;
        RECT 35.225 -115.030 35.605 -114.650 ;
        RECT 39.225 -114.695 39.605 -114.650 ;
        RECT 44.725 -114.695 45.105 -114.650 ;
        RECT 39.175 -115.010 45.110 -114.695 ;
        RECT 39.225 -115.030 39.605 -115.010 ;
        RECT 44.725 -115.030 45.105 -115.010 ;
        RECT 48.725 -115.030 49.105 -114.650 ;
        RECT 52.725 -115.030 53.105 -114.650 ;
        RECT 69.845 -115.010 70.225 -114.630 ;
        RECT 73.845 -115.010 74.225 -114.630 ;
        RECT 77.845 -114.675 78.225 -114.630 ;
        RECT 83.345 -114.675 83.725 -114.630 ;
        RECT 77.795 -114.990 83.730 -114.675 ;
        RECT 77.845 -115.010 78.225 -114.990 ;
        RECT 83.345 -115.010 83.725 -114.990 ;
        RECT 87.345 -115.010 87.725 -114.630 ;
        RECT 91.345 -115.010 91.725 -114.630 ;
        RECT 97.055 -114.710 98.795 -114.420 ;
        RECT 100.845 -114.760 102.045 -114.470 ;
        RECT 103.555 -114.800 106.185 -114.345 ;
        RECT 107.765 -114.695 108.145 -114.315 ;
        RECT 61.935 -115.635 82.710 -115.260 ;
        RECT 32.450 -116.245 59.760 -115.905 ;
        RECT 12.065 -116.950 19.325 -116.650 ;
        RECT 12.620 -117.485 16.705 -117.215 ;
        RECT 23.025 -117.250 26.775 -116.975 ;
        RECT 60.965 -116.990 92.930 -116.600 ;
        RECT 105.740 -117.230 108.870 -116.955 ;
        RECT 109.615 -116.990 109.995 -109.830 ;
        RECT 110.855 -112.290 117.595 -111.990 ;
        RECT 111.445 -114.085 114.900 -113.645 ;
        RECT 117.905 -114.245 118.285 -113.865 ;
        RECT 116.305 -114.760 117.505 -114.470 ;
        RECT 123.225 -114.695 123.605 -114.315 ;
        RECT 110.260 -115.470 126.180 -115.170 ;
        RECT 110.795 -116.215 127.740 -115.915 ;
        RECT 57.810 -117.355 85.370 -117.345 ;
        RECT 28.080 -117.375 46.750 -117.365 ;
        RECT 57.810 -117.375 94.375 -117.355 ;
        RECT 28.080 -117.665 94.375 -117.375 ;
        RECT 28.080 -117.685 58.100 -117.665 ;
        RECT 111.990 -118.125 116.120 -117.825 ;
        RECT -4.020 -123.975 -3.640 -118.145 ;
        RECT 0.235 -119.325 10.890 -118.990 ;
        RECT 0.205 -120.645 1.985 -120.355 ;
        RECT 7.580 -120.675 8.890 -120.355 ;
        RECT -1.065 -121.260 -0.685 -120.880 ;
        RECT 5.390 -121.230 5.770 -120.850 ;
        RECT -3.270 -123.975 0.825 -123.970 ;
        RECT 11.440 -123.975 11.820 -118.145 ;
        RECT 63.030 -118.355 94.775 -118.335 ;
        RECT 16.280 -118.745 22.670 -118.455 ;
        RECT 27.550 -118.605 94.775 -118.355 ;
        RECT 27.550 -118.625 63.460 -118.605 ;
        RECT 98.995 -118.725 105.385 -118.435 ;
        RECT 15.695 -119.325 26.200 -118.990 ;
        RECT 51.170 -119.190 61.720 -118.855 ;
        RECT 98.410 -119.305 108.890 -118.970 ;
        RECT 31.765 -119.830 35.065 -119.450 ;
        RECT 35.765 -119.830 39.065 -119.450 ;
        RECT 45.265 -119.830 48.565 -119.450 ;
        RECT 49.265 -119.830 52.565 -119.450 ;
        RECT 68.380 -119.810 69.685 -119.430 ;
        RECT 74.385 -119.810 77.685 -119.430 ;
        RECT 78.385 -119.810 79.745 -119.430 ;
        RECT 81.720 -119.810 83.185 -119.430 ;
        RECT 83.885 -119.810 87.185 -119.430 ;
        RECT 91.885 -119.810 93.065 -119.430 ;
        RECT 31.225 -120.175 31.605 -120.140 ;
        RECT 13.260 -120.660 13.640 -120.280 ;
        RECT 15.665 -120.645 17.445 -120.355 ;
        RECT 18.920 -120.555 20.110 -120.270 ;
        RECT 23.040 -120.675 24.350 -120.355 ;
        RECT 30.960 -120.485 33.970 -120.175 ;
        RECT 31.225 -120.520 31.605 -120.485 ;
        RECT 35.225 -120.520 36.315 -120.140 ;
        RECT 39.225 -120.145 39.605 -120.140 ;
        RECT 36.745 -120.510 39.610 -120.145 ;
        RECT 44.725 -120.165 45.105 -120.140 ;
        RECT 44.710 -120.485 46.855 -120.165 ;
        RECT 39.225 -120.520 39.605 -120.510 ;
        RECT 44.725 -120.520 45.105 -120.485 ;
        RECT 47.770 -120.520 49.105 -120.140 ;
        RECT 52.725 -120.160 53.105 -120.140 ;
        RECT 69.845 -120.155 70.225 -120.120 ;
        RECT 50.260 -120.480 53.170 -120.160 ;
        RECT 69.580 -120.465 72.590 -120.155 ;
        RECT 52.725 -120.520 53.105 -120.480 ;
        RECT 69.845 -120.500 70.225 -120.465 ;
        RECT 73.845 -120.500 74.935 -120.120 ;
        RECT 77.845 -120.125 78.225 -120.120 ;
        RECT 75.365 -120.490 78.230 -120.125 ;
        RECT 83.345 -120.145 83.725 -120.120 ;
        RECT 83.330 -120.465 85.475 -120.145 ;
        RECT 77.845 -120.500 78.225 -120.490 ;
        RECT 83.345 -120.500 83.725 -120.465 ;
        RECT 86.390 -120.500 87.725 -120.120 ;
        RECT 91.345 -120.140 91.725 -120.120 ;
        RECT 88.880 -120.460 91.790 -120.140 ;
        RECT 91.345 -120.500 91.725 -120.460 ;
        RECT 95.975 -120.640 96.355 -120.260 ;
        RECT 98.380 -120.625 100.160 -120.335 ;
        RECT 101.635 -120.535 102.825 -120.250 ;
        RECT 105.755 -120.655 107.065 -120.335 ;
        RECT 14.395 -121.260 14.775 -120.880 ;
        RECT 18.140 -121.220 18.520 -120.840 ;
        RECT 20.850 -121.230 21.230 -120.850 ;
        RECT 22.260 -121.385 25.440 -121.065 ;
        RECT 97.110 -121.240 97.490 -120.860 ;
        RECT 100.855 -121.200 101.235 -120.820 ;
        RECT 103.565 -121.210 103.945 -120.830 ;
        RECT 104.975 -121.365 108.155 -121.045 ;
        RECT 31.765 -121.830 33.050 -121.450 ;
        RECT 51.080 -121.830 52.565 -121.450 ;
        RECT 68.195 -121.810 69.685 -121.430 ;
        RECT 91.885 -121.810 92.960 -121.430 ;
        RECT 31.225 -122.520 32.315 -122.140 ;
        RECT 33.270 -122.510 34.790 -122.150 ;
        RECT 35.710 -122.515 48.560 -122.180 ;
        RECT 52.725 -122.185 53.105 -122.140 ;
        RECT 51.990 -122.485 53.300 -122.185 ;
        RECT 52.725 -122.520 53.105 -122.485 ;
        RECT 69.845 -122.500 70.935 -122.120 ;
        RECT 71.890 -122.490 73.410 -122.130 ;
        RECT 74.330 -122.495 87.180 -122.160 ;
        RECT 91.345 -122.165 91.725 -122.120 ;
        RECT 90.610 -122.465 91.920 -122.165 ;
        RECT 91.345 -122.500 91.725 -122.465 ;
        RECT 60.405 -123.030 93.355 -122.995 ;
        RECT 28.080 -123.360 93.355 -123.030 ;
        RECT 28.080 -123.380 61.160 -123.360 ;
        RECT 95.150 -123.370 99.410 -123.015 ;
        RECT 93.355 -123.955 99.000 -123.950 ;
        RECT 109.615 -123.955 109.995 -118.125 ;
        RECT 118.495 -118.175 122.995 -117.865 ;
        RECT 114.455 -118.725 120.845 -118.435 ;
        RECT 113.220 -119.890 116.140 -119.590 ;
        RECT 119.685 -119.905 123.055 -119.605 ;
        RECT 111.435 -120.640 111.815 -120.260 ;
        RECT 117.095 -120.535 118.285 -120.250 ;
        RECT 116.315 -121.200 116.695 -120.820 ;
        RECT 120.435 -121.365 123.615 -121.045 ;
        RECT 110.715 -122.450 114.865 -122.180 ;
        RECT 110.365 -123.955 114.460 -123.950 ;
        RECT 66.700 -123.960 99.000 -123.955 ;
        RECT 109.245 -123.960 114.460 -123.955 ;
        RECT 12.190 -123.975 16.285 -123.970 ;
        RECT 66.700 -123.975 124.275 -123.960 ;
        RECT -4.390 -123.980 0.825 -123.975 ;
        RECT 11.070 -123.980 16.285 -123.975 ;
        RECT 26.530 -123.980 124.275 -123.975 ;
        RECT -4.390 -124.855 124.275 -123.980 ;
        RECT -4.390 -124.875 66.780 -124.855 ;
        RECT -4.440 -128.900 67.950 -128.760 ;
        RECT -4.440 -129.660 124.275 -128.900 ;
        RECT -4.070 -136.820 -3.690 -129.660 ;
        RECT 1.505 -134.115 1.885 -133.735 ;
        RECT 8.405 -134.125 8.785 -133.745 ;
        RECT -1.170 -134.540 0.570 -134.250 ;
        RECT 5.330 -134.620 7.940 -134.195 ;
        RECT 7.515 -137.060 10.620 -136.785 ;
        RECT 11.390 -136.820 11.770 -129.660 ;
        RECT 67.920 -129.800 124.275 -129.660 ;
        RECT 28.030 -130.785 65.580 -130.645 ;
        RECT 28.030 -130.930 93.680 -130.785 ;
        RECT 64.905 -131.070 93.680 -130.930 ;
        RECT 95.350 -131.090 102.055 -130.790 ;
        RECT 31.735 -131.840 32.935 -131.460 ;
        RECT 34.690 -132.055 36.965 -131.545 ;
        RECT 39.590 -132.055 41.890 -131.545 ;
        RECT 44.185 -132.055 46.465 -131.545 ;
        RECT 51.260 -131.740 52.495 -131.360 ;
        RECT 68.210 -131.980 69.665 -131.600 ;
        RECT 52.675 -132.095 53.055 -132.060 ;
        RECT 31.175 -132.200 31.555 -132.160 ;
        RECT 31.105 -132.505 33.940 -132.200 ;
        RECT 49.920 -132.405 53.055 -132.095 ;
        RECT 73.360 -132.195 75.635 -131.685 ;
        RECT 78.260 -132.195 80.560 -131.685 ;
        RECT 82.855 -132.195 85.135 -131.685 ;
        RECT 91.905 -131.880 93.185 -131.500 ;
        RECT 91.345 -132.235 91.725 -132.200 ;
        RECT 69.845 -132.340 70.225 -132.300 ;
        RECT 52.675 -132.440 53.055 -132.405 ;
        RECT 31.175 -132.540 31.555 -132.505 ;
        RECT 69.775 -132.645 72.610 -132.340 ;
        RECT 88.590 -132.545 91.725 -132.235 ;
        RECT 91.345 -132.580 91.725 -132.545 ;
        RECT 69.845 -132.680 70.225 -132.645 ;
        RECT 13.220 -133.915 16.625 -133.475 ;
        RECT 16.965 -134.115 17.345 -133.735 ;
        RECT 19.680 -134.075 20.060 -133.695 ;
        RECT 23.865 -134.125 24.245 -133.745 ;
        RECT 31.735 -134.140 34.995 -133.760 ;
        RECT 35.735 -134.140 38.995 -133.760 ;
        RECT 45.235 -134.140 48.495 -133.760 ;
        RECT 49.235 -134.140 52.495 -133.760 ;
        RECT 14.290 -134.540 16.030 -134.250 ;
        RECT 18.080 -134.590 19.280 -134.300 ;
        RECT 20.790 -134.620 23.385 -134.245 ;
        RECT 25.000 -134.525 25.380 -134.145 ;
        RECT 68.370 -134.280 69.665 -133.900 ;
        RECT 74.405 -134.280 77.665 -133.900 ;
        RECT 78.405 -134.280 79.590 -133.900 ;
        RECT 81.855 -134.280 83.165 -133.900 ;
        RECT 83.905 -134.280 87.165 -133.900 ;
        RECT 91.905 -134.280 92.920 -133.900 ;
        RECT 95.985 -134.035 99.400 -133.615 ;
        RECT 99.730 -134.255 100.110 -133.875 ;
        RECT 102.445 -134.215 102.825 -133.835 ;
        RECT 106.630 -134.265 107.010 -133.885 ;
        RECT 31.175 -134.840 31.555 -134.460 ;
        RECT 35.175 -134.840 35.555 -134.460 ;
        RECT 39.175 -134.505 39.555 -134.460 ;
        RECT 44.675 -134.505 45.055 -134.460 ;
        RECT 39.125 -134.820 45.060 -134.505 ;
        RECT 39.175 -134.840 39.555 -134.820 ;
        RECT 44.675 -134.840 45.055 -134.820 ;
        RECT 48.675 -134.840 49.055 -134.460 ;
        RECT 52.675 -134.840 53.055 -134.460 ;
        RECT 69.845 -134.980 70.225 -134.600 ;
        RECT 73.845 -134.980 74.225 -134.600 ;
        RECT 77.845 -134.645 78.225 -134.600 ;
        RECT 83.345 -134.645 83.725 -134.600 ;
        RECT 77.795 -134.960 83.730 -134.645 ;
        RECT 77.845 -134.980 78.225 -134.960 ;
        RECT 83.345 -134.980 83.725 -134.960 ;
        RECT 87.345 -134.980 87.725 -134.600 ;
        RECT 91.345 -134.980 91.725 -134.600 ;
        RECT 97.055 -134.680 98.795 -134.390 ;
        RECT 100.845 -134.730 102.045 -134.440 ;
        RECT 103.555 -134.770 106.185 -134.315 ;
        RECT 107.765 -134.665 108.145 -134.285 ;
        RECT 61.935 -135.605 82.710 -135.230 ;
        RECT 32.400 -136.055 59.710 -135.715 ;
        RECT 12.015 -136.760 19.275 -136.460 ;
        RECT 12.570 -137.295 16.655 -137.025 ;
        RECT 22.975 -137.060 26.725 -136.785 ;
        RECT 60.965 -136.960 92.930 -136.570 ;
        RECT 28.030 -137.185 46.700 -137.175 ;
        RECT 28.030 -137.315 58.050 -137.185 ;
        RECT 105.740 -137.200 108.870 -136.925 ;
        RECT 109.615 -136.960 109.995 -129.800 ;
        RECT 110.855 -132.260 117.595 -131.960 ;
        RECT 111.445 -134.055 114.900 -133.615 ;
        RECT 117.905 -134.215 118.285 -133.835 ;
        RECT 116.305 -134.730 117.505 -134.440 ;
        RECT 123.225 -134.665 123.605 -134.285 ;
        RECT 110.260 -135.440 126.180 -135.140 ;
        RECT 110.795 -136.185 127.740 -135.885 ;
        RECT 28.030 -137.325 85.370 -137.315 ;
        RECT 28.030 -137.495 94.375 -137.325 ;
        RECT 57.810 -137.635 94.375 -137.495 ;
        RECT -4.070 -143.785 -3.690 -137.955 ;
        RECT 0.185 -139.135 10.840 -138.800 ;
        RECT 0.155 -140.455 1.935 -140.165 ;
        RECT 7.530 -140.485 8.840 -140.165 ;
        RECT -1.115 -141.070 -0.735 -140.690 ;
        RECT 5.340 -141.040 5.720 -140.660 ;
        RECT -3.320 -143.785 0.775 -143.780 ;
        RECT 11.390 -143.785 11.770 -137.955 ;
        RECT 111.990 -138.095 116.120 -137.795 ;
        RECT 16.230 -138.555 22.620 -138.265 ;
        RECT 27.500 -138.305 63.410 -138.165 ;
        RECT 27.500 -138.435 94.775 -138.305 ;
        RECT 63.030 -138.575 94.775 -138.435 ;
        RECT 15.645 -139.135 26.150 -138.800 ;
        RECT 51.120 -139.000 61.670 -138.665 ;
        RECT 98.995 -138.695 105.385 -138.405 ;
        RECT 31.715 -139.640 35.015 -139.260 ;
        RECT 35.715 -139.640 39.015 -139.260 ;
        RECT 45.215 -139.640 48.515 -139.260 ;
        RECT 49.215 -139.640 52.515 -139.260 ;
        RECT 98.410 -139.275 108.890 -138.940 ;
        RECT 68.380 -139.780 69.685 -139.400 ;
        RECT 74.385 -139.780 77.685 -139.400 ;
        RECT 78.385 -139.780 79.745 -139.400 ;
        RECT 81.720 -139.780 83.185 -139.400 ;
        RECT 83.885 -139.780 87.185 -139.400 ;
        RECT 91.885 -139.780 93.065 -139.400 ;
        RECT 31.175 -139.985 31.555 -139.950 ;
        RECT 13.210 -140.470 13.590 -140.090 ;
        RECT 15.615 -140.455 17.395 -140.165 ;
        RECT 18.870 -140.365 20.060 -140.080 ;
        RECT 22.990 -140.485 24.300 -140.165 ;
        RECT 30.910 -140.295 33.920 -139.985 ;
        RECT 31.175 -140.330 31.555 -140.295 ;
        RECT 35.175 -140.330 36.265 -139.950 ;
        RECT 39.175 -139.955 39.555 -139.950 ;
        RECT 36.695 -140.320 39.560 -139.955 ;
        RECT 44.675 -139.975 45.055 -139.950 ;
        RECT 44.660 -140.295 46.805 -139.975 ;
        RECT 39.175 -140.330 39.555 -140.320 ;
        RECT 44.675 -140.330 45.055 -140.295 ;
        RECT 47.720 -140.330 49.055 -139.950 ;
        RECT 52.675 -139.970 53.055 -139.950 ;
        RECT 50.210 -140.290 53.120 -139.970 ;
        RECT 69.845 -140.125 70.225 -140.090 ;
        RECT 52.675 -140.330 53.055 -140.290 ;
        RECT 69.580 -140.435 72.590 -140.125 ;
        RECT 69.845 -140.470 70.225 -140.435 ;
        RECT 73.845 -140.470 74.935 -140.090 ;
        RECT 77.845 -140.095 78.225 -140.090 ;
        RECT 75.365 -140.460 78.230 -140.095 ;
        RECT 83.345 -140.115 83.725 -140.090 ;
        RECT 83.330 -140.435 85.475 -140.115 ;
        RECT 77.845 -140.470 78.225 -140.460 ;
        RECT 83.345 -140.470 83.725 -140.435 ;
        RECT 86.390 -140.470 87.725 -140.090 ;
        RECT 91.345 -140.110 91.725 -140.090 ;
        RECT 88.880 -140.430 91.790 -140.110 ;
        RECT 91.345 -140.470 91.725 -140.430 ;
        RECT 95.975 -140.610 96.355 -140.230 ;
        RECT 98.380 -140.595 100.160 -140.305 ;
        RECT 101.635 -140.505 102.825 -140.220 ;
        RECT 105.755 -140.625 107.065 -140.305 ;
        RECT 14.345 -141.070 14.725 -140.690 ;
        RECT 18.090 -141.030 18.470 -140.650 ;
        RECT 20.800 -141.040 21.180 -140.660 ;
        RECT 22.210 -141.195 25.390 -140.875 ;
        RECT 97.110 -141.210 97.490 -140.830 ;
        RECT 100.855 -141.170 101.235 -140.790 ;
        RECT 103.565 -141.180 103.945 -140.800 ;
        RECT 31.715 -141.640 33.000 -141.260 ;
        RECT 51.030 -141.640 52.515 -141.260 ;
        RECT 104.975 -141.335 108.155 -141.015 ;
        RECT 68.195 -141.780 69.685 -141.400 ;
        RECT 91.885 -141.780 92.960 -141.400 ;
        RECT 31.175 -142.330 32.265 -141.950 ;
        RECT 33.220 -142.320 34.740 -141.960 ;
        RECT 35.660 -142.325 48.510 -141.990 ;
        RECT 52.675 -141.995 53.055 -141.950 ;
        RECT 51.940 -142.295 53.250 -141.995 ;
        RECT 52.675 -142.330 53.055 -142.295 ;
        RECT 69.845 -142.470 70.935 -142.090 ;
        RECT 71.890 -142.460 73.410 -142.100 ;
        RECT 74.330 -142.465 87.180 -142.130 ;
        RECT 91.345 -142.135 91.725 -142.090 ;
        RECT 90.610 -142.435 91.920 -142.135 ;
        RECT 91.345 -142.470 91.725 -142.435 ;
        RECT 28.030 -142.965 61.110 -142.840 ;
        RECT 28.030 -143.190 93.355 -142.965 ;
        RECT 60.405 -143.330 93.355 -143.190 ;
        RECT 95.150 -143.340 99.410 -142.985 ;
        RECT 12.140 -143.785 16.235 -143.780 ;
        RECT -4.440 -143.790 0.775 -143.785 ;
        RECT 11.020 -143.790 16.235 -143.785 ;
        RECT 26.480 -143.790 66.730 -143.785 ;
        RECT -4.440 -143.925 66.730 -143.790 ;
        RECT 93.355 -143.925 99.000 -143.920 ;
        RECT 109.615 -143.925 109.995 -138.095 ;
        RECT 118.495 -138.145 122.995 -137.835 ;
        RECT 114.455 -138.695 120.845 -138.405 ;
        RECT 113.220 -139.860 116.140 -139.560 ;
        RECT 119.685 -139.875 123.055 -139.575 ;
        RECT 111.435 -140.610 111.815 -140.230 ;
        RECT 117.095 -140.505 118.285 -140.220 ;
        RECT 116.315 -141.170 116.695 -140.790 ;
        RECT 120.435 -141.335 123.615 -141.015 ;
        RECT 110.715 -142.420 114.865 -142.150 ;
        RECT 110.365 -143.925 114.460 -143.920 ;
        RECT -4.440 -143.930 99.000 -143.925 ;
        RECT 109.245 -143.930 114.460 -143.925 ;
        RECT -4.440 -144.685 124.275 -143.930 ;
        RECT 66.700 -144.825 124.275 -144.685 ;
        RECT -4.470 -148.565 67.920 -148.555 ;
        RECT -4.470 -149.455 124.275 -148.565 ;
        RECT -4.100 -156.615 -3.720 -149.455 ;
        RECT 1.475 -153.910 1.855 -153.530 ;
        RECT 8.375 -153.920 8.755 -153.540 ;
        RECT -1.200 -154.335 0.540 -154.045 ;
        RECT 5.300 -154.415 7.910 -153.990 ;
        RECT 7.485 -156.855 10.590 -156.580 ;
        RECT 11.360 -156.615 11.740 -149.455 ;
        RECT 67.920 -149.465 124.275 -149.455 ;
        RECT 28.000 -150.450 65.550 -150.440 ;
        RECT 28.000 -150.725 93.680 -150.450 ;
        RECT 64.905 -150.735 93.680 -150.725 ;
        RECT 95.350 -150.755 102.055 -150.455 ;
        RECT 31.705 -151.635 32.905 -151.255 ;
        RECT 34.660 -151.850 36.935 -151.340 ;
        RECT 39.560 -151.850 41.860 -151.340 ;
        RECT 44.155 -151.850 46.435 -151.340 ;
        RECT 51.230 -151.535 52.465 -151.155 ;
        RECT 68.210 -151.645 69.665 -151.265 ;
        RECT 52.645 -151.890 53.025 -151.855 ;
        RECT 73.360 -151.860 75.635 -151.350 ;
        RECT 78.260 -151.860 80.560 -151.350 ;
        RECT 82.855 -151.860 85.135 -151.350 ;
        RECT 91.905 -151.545 93.185 -151.165 ;
        RECT 31.145 -151.995 31.525 -151.955 ;
        RECT 31.075 -152.300 33.910 -151.995 ;
        RECT 49.890 -152.200 53.025 -151.890 ;
        RECT 91.345 -151.900 91.725 -151.865 ;
        RECT 69.845 -152.005 70.225 -151.965 ;
        RECT 52.645 -152.235 53.025 -152.200 ;
        RECT 31.145 -152.335 31.525 -152.300 ;
        RECT 69.775 -152.310 72.610 -152.005 ;
        RECT 88.590 -152.210 91.725 -151.900 ;
        RECT 91.345 -152.245 91.725 -152.210 ;
        RECT 69.845 -152.345 70.225 -152.310 ;
        RECT 13.190 -153.710 16.595 -153.270 ;
        RECT 16.935 -153.910 17.315 -153.530 ;
        RECT 19.650 -153.870 20.030 -153.490 ;
        RECT 23.835 -153.920 24.215 -153.540 ;
        RECT 31.705 -153.935 34.965 -153.555 ;
        RECT 35.705 -153.935 38.965 -153.555 ;
        RECT 45.205 -153.935 48.465 -153.555 ;
        RECT 49.205 -153.935 52.465 -153.555 ;
        RECT 14.260 -154.335 16.000 -154.045 ;
        RECT 18.050 -154.385 19.250 -154.095 ;
        RECT 20.760 -154.415 23.355 -154.040 ;
        RECT 24.970 -154.320 25.350 -153.940 ;
        RECT 68.370 -153.945 69.665 -153.565 ;
        RECT 74.405 -153.945 77.665 -153.565 ;
        RECT 78.405 -153.945 79.590 -153.565 ;
        RECT 81.855 -153.945 83.165 -153.565 ;
        RECT 83.905 -153.945 87.165 -153.565 ;
        RECT 91.905 -153.945 92.920 -153.565 ;
        RECT 95.985 -153.700 99.400 -153.280 ;
        RECT 99.730 -153.920 100.110 -153.540 ;
        RECT 102.445 -153.880 102.825 -153.500 ;
        RECT 106.630 -153.930 107.010 -153.550 ;
        RECT 31.145 -154.635 31.525 -154.255 ;
        RECT 35.145 -154.635 35.525 -154.255 ;
        RECT 39.145 -154.300 39.525 -154.255 ;
        RECT 44.645 -154.300 45.025 -154.255 ;
        RECT 39.095 -154.615 45.030 -154.300 ;
        RECT 39.145 -154.635 39.525 -154.615 ;
        RECT 44.645 -154.635 45.025 -154.615 ;
        RECT 48.645 -154.635 49.025 -154.255 ;
        RECT 52.645 -154.635 53.025 -154.255 ;
        RECT 69.845 -154.645 70.225 -154.265 ;
        RECT 73.845 -154.645 74.225 -154.265 ;
        RECT 77.845 -154.310 78.225 -154.265 ;
        RECT 83.345 -154.310 83.725 -154.265 ;
        RECT 77.795 -154.625 83.730 -154.310 ;
        RECT 77.845 -154.645 78.225 -154.625 ;
        RECT 83.345 -154.645 83.725 -154.625 ;
        RECT 87.345 -154.645 87.725 -154.265 ;
        RECT 91.345 -154.645 91.725 -154.265 ;
        RECT 97.055 -154.345 98.795 -154.055 ;
        RECT 100.845 -154.395 102.045 -154.105 ;
        RECT 103.555 -154.435 106.185 -153.980 ;
        RECT 107.765 -154.330 108.145 -153.950 ;
        RECT 61.935 -155.270 82.710 -154.895 ;
        RECT 32.370 -155.850 59.680 -155.510 ;
        RECT 11.985 -156.555 19.245 -156.255 ;
        RECT 12.540 -157.090 16.625 -156.820 ;
        RECT 22.945 -156.855 26.695 -156.580 ;
        RECT 60.965 -156.625 92.930 -156.235 ;
        RECT 105.740 -156.865 108.870 -156.590 ;
        RECT 109.615 -156.625 109.995 -149.465 ;
        RECT 110.855 -151.925 117.595 -151.625 ;
        RECT 111.445 -153.720 114.900 -153.280 ;
        RECT 117.905 -153.880 118.285 -153.500 ;
        RECT 116.305 -154.395 117.505 -154.105 ;
        RECT 123.225 -154.330 123.605 -153.950 ;
        RECT 110.260 -155.105 126.180 -154.805 ;
        RECT 110.795 -155.850 127.740 -155.550 ;
        RECT 28.000 -156.980 46.670 -156.970 ;
        RECT 28.000 -156.990 85.370 -156.980 ;
        RECT 28.000 -157.290 94.375 -156.990 ;
        RECT 57.810 -157.300 94.375 -157.290 ;
        RECT -4.100 -163.580 -3.720 -157.750 ;
        RECT 0.155 -158.930 10.810 -158.595 ;
        RECT 0.125 -160.250 1.905 -159.960 ;
        RECT 7.500 -160.280 8.810 -159.960 ;
        RECT -1.145 -160.865 -0.765 -160.485 ;
        RECT 5.310 -160.835 5.690 -160.455 ;
        RECT -3.350 -163.580 0.745 -163.575 ;
        RECT 11.360 -163.580 11.740 -157.750 ;
        RECT 111.990 -157.760 116.120 -157.460 ;
        RECT 27.470 -157.970 63.380 -157.960 ;
        RECT 16.200 -158.350 22.590 -158.060 ;
        RECT 27.470 -158.230 94.775 -157.970 ;
        RECT 63.030 -158.240 94.775 -158.230 ;
        RECT 98.995 -158.360 105.385 -158.070 ;
        RECT 15.615 -158.930 26.120 -158.595 ;
        RECT 51.090 -158.795 61.640 -158.460 ;
        RECT 98.410 -158.940 108.890 -158.605 ;
        RECT 31.685 -159.435 34.985 -159.055 ;
        RECT 35.685 -159.435 38.985 -159.055 ;
        RECT 45.185 -159.435 48.485 -159.055 ;
        RECT 49.185 -159.435 52.485 -159.055 ;
        RECT 68.380 -159.445 69.685 -159.065 ;
        RECT 74.385 -159.445 77.685 -159.065 ;
        RECT 78.385 -159.445 79.745 -159.065 ;
        RECT 81.720 -159.445 83.185 -159.065 ;
        RECT 83.885 -159.445 87.185 -159.065 ;
        RECT 91.885 -159.445 93.065 -159.065 ;
        RECT 31.145 -159.780 31.525 -159.745 ;
        RECT 13.180 -160.265 13.560 -159.885 ;
        RECT 15.585 -160.250 17.365 -159.960 ;
        RECT 18.840 -160.160 20.030 -159.875 ;
        RECT 22.960 -160.280 24.270 -159.960 ;
        RECT 30.880 -160.090 33.890 -159.780 ;
        RECT 31.145 -160.125 31.525 -160.090 ;
        RECT 35.145 -160.125 36.235 -159.745 ;
        RECT 39.145 -159.750 39.525 -159.745 ;
        RECT 36.665 -160.115 39.530 -159.750 ;
        RECT 44.645 -159.770 45.025 -159.745 ;
        RECT 44.630 -160.090 46.775 -159.770 ;
        RECT 39.145 -160.125 39.525 -160.115 ;
        RECT 44.645 -160.125 45.025 -160.090 ;
        RECT 47.690 -160.125 49.025 -159.745 ;
        RECT 52.645 -159.765 53.025 -159.745 ;
        RECT 50.180 -160.085 53.090 -159.765 ;
        RECT 69.845 -159.790 70.225 -159.755 ;
        RECT 52.645 -160.125 53.025 -160.085 ;
        RECT 69.580 -160.100 72.590 -159.790 ;
        RECT 69.845 -160.135 70.225 -160.100 ;
        RECT 73.845 -160.135 74.935 -159.755 ;
        RECT 77.845 -159.760 78.225 -159.755 ;
        RECT 75.365 -160.125 78.230 -159.760 ;
        RECT 83.345 -159.780 83.725 -159.755 ;
        RECT 83.330 -160.100 85.475 -159.780 ;
        RECT 77.845 -160.135 78.225 -160.125 ;
        RECT 83.345 -160.135 83.725 -160.100 ;
        RECT 86.390 -160.135 87.725 -159.755 ;
        RECT 91.345 -159.775 91.725 -159.755 ;
        RECT 88.880 -160.095 91.790 -159.775 ;
        RECT 91.345 -160.135 91.725 -160.095 ;
        RECT 95.975 -160.275 96.355 -159.895 ;
        RECT 98.380 -160.260 100.160 -159.970 ;
        RECT 101.635 -160.170 102.825 -159.885 ;
        RECT 105.755 -160.290 107.065 -159.970 ;
        RECT 14.315 -160.865 14.695 -160.485 ;
        RECT 18.060 -160.825 18.440 -160.445 ;
        RECT 20.770 -160.835 21.150 -160.455 ;
        RECT 22.180 -160.990 25.360 -160.670 ;
        RECT 97.110 -160.875 97.490 -160.495 ;
        RECT 100.855 -160.835 101.235 -160.455 ;
        RECT 103.565 -160.845 103.945 -160.465 ;
        RECT 104.975 -161.000 108.155 -160.680 ;
        RECT 31.685 -161.435 32.970 -161.055 ;
        RECT 51.000 -161.435 52.485 -161.055 ;
        RECT 68.195 -161.445 69.685 -161.065 ;
        RECT 91.885 -161.445 92.960 -161.065 ;
        RECT 31.145 -162.125 32.235 -161.745 ;
        RECT 33.190 -162.115 34.710 -161.755 ;
        RECT 35.630 -162.120 48.480 -161.785 ;
        RECT 52.645 -161.790 53.025 -161.745 ;
        RECT 51.910 -162.090 53.220 -161.790 ;
        RECT 52.645 -162.125 53.025 -162.090 ;
        RECT 69.845 -162.135 70.935 -161.755 ;
        RECT 71.890 -162.125 73.410 -161.765 ;
        RECT 74.330 -162.130 87.180 -161.795 ;
        RECT 91.345 -161.800 91.725 -161.755 ;
        RECT 90.610 -162.100 91.920 -161.800 ;
        RECT 91.345 -162.135 91.725 -162.100 ;
        RECT 60.405 -162.635 93.355 -162.630 ;
        RECT 28.000 -162.985 93.355 -162.635 ;
        RECT 60.405 -162.995 93.355 -162.985 ;
        RECT 95.150 -163.005 99.410 -162.650 ;
        RECT 12.110 -163.580 16.205 -163.575 ;
        RECT -4.470 -163.585 0.745 -163.580 ;
        RECT 10.990 -163.585 16.205 -163.580 ;
        RECT 26.450 -163.585 66.700 -163.580 ;
        RECT -4.470 -163.590 66.700 -163.585 ;
        RECT 93.355 -163.590 99.000 -163.585 ;
        RECT 109.615 -163.590 109.995 -157.760 ;
        RECT 118.495 -157.810 122.995 -157.500 ;
        RECT 114.455 -158.360 120.845 -158.070 ;
        RECT 113.220 -159.525 116.140 -159.225 ;
        RECT 119.685 -159.540 123.055 -159.240 ;
        RECT 111.435 -160.275 111.815 -159.895 ;
        RECT 117.095 -160.170 118.285 -159.885 ;
        RECT 116.315 -160.835 116.695 -160.455 ;
        RECT 120.435 -161.000 123.615 -160.680 ;
        RECT 110.715 -162.085 114.865 -161.815 ;
        RECT 110.365 -163.590 114.460 -163.585 ;
        RECT -4.470 -163.595 99.000 -163.590 ;
        RECT 109.245 -163.595 114.460 -163.590 ;
        RECT -4.470 -164.480 124.275 -163.595 ;
        RECT 66.700 -164.490 124.275 -164.480 ;
        RECT 67.365 -173.450 70.765 -173.015 ;
        RECT 73.825 -173.615 74.205 -173.235 ;
        RECT 72.225 -174.130 73.425 -173.840 ;
        RECT 79.145 -174.065 79.525 -173.685 ;
        RECT 62.870 -174.840 80.195 -174.540 ;
        RECT 62.630 -175.585 80.195 -175.285 ;
        RECT 64.490 -176.300 73.420 -176.000 ;
        RECT 64.460 -176.835 70.800 -176.565 ;
        RECT 67.910 -177.495 72.040 -177.195 ;
        RECT 74.415 -177.545 78.915 -177.235 ;
        RECT 70.375 -178.095 76.765 -177.805 ;
        RECT 69.140 -179.260 72.060 -178.960 ;
        RECT 75.605 -179.275 78.975 -178.975 ;
        RECT 67.355 -180.010 67.735 -179.630 ;
        RECT 73.015 -179.905 74.205 -179.620 ;
        RECT 72.235 -180.570 72.615 -180.190 ;
        RECT 76.355 -180.735 79.535 -180.415 ;
      LAYER Metal2 ;
        RECT -1.005 135.500 -0.705 142.430 ;
        RECT 0.305 136.100 0.605 142.450 ;
        RECT 1.620 136.130 1.915 142.955 ;
        RECT 5.460 135.500 5.760 142.440 ;
        RECT 7.670 136.075 7.975 142.435 ;
        RECT 8.520 136.075 8.820 142.895 ;
        RECT 10.330 139.520 10.710 139.900 ;
        RECT 12.115 138.100 12.435 140.230 ;
        RECT 10.545 134.810 10.925 137.830 ;
        RECT 12.725 137.260 13.005 139.665 ;
        RECT 13.335 136.105 13.635 143.145 ;
        RECT 14.455 135.500 14.755 142.430 ;
        RECT 15.765 136.100 16.065 142.450 ;
        RECT 16.360 137.975 16.685 143.135 ;
        RECT 17.080 136.130 17.375 142.955 ;
        RECT 18.210 135.590 18.510 142.400 ;
        RECT 19.000 136.185 19.310 142.375 ;
        RECT 19.795 136.115 20.095 142.945 ;
        RECT 20.920 135.500 21.220 142.440 ;
        RECT 22.370 135.375 22.650 138.410 ;
        RECT 23.130 136.075 23.450 142.435 ;
        RECT 23.980 136.075 24.280 142.895 ;
        RECT 25.120 135.330 25.420 142.485 ;
        RECT 25.755 137.475 26.135 137.855 ;
        RECT 26.460 133.360 26.820 139.920 ;
        RECT 27.600 138.110 27.925 139.975 ;
        RECT 28.265 134.765 28.725 139.450 ;
        RECT 29.050 137.310 29.500 146.130 ;
        RECT 31.235 139.135 31.665 142.125 ;
        RECT 28.980 133.420 29.360 133.800 ;
        RECT 31.870 133.440 32.250 134.815 ;
        RECT 32.640 134.260 32.955 145.310 ;
        RECT 33.655 144.005 33.945 146.065 ;
        RECT 36.440 144.605 36.915 147.655 ;
        RECT 41.395 144.515 41.805 147.610 ;
        RECT 33.575 136.150 33.900 138.520 ;
        RECT 35.225 138.195 35.625 142.160 ;
        RECT 34.310 132.410 34.655 134.870 ;
        RECT 35.945 134.090 36.270 136.855 ;
        RECT 36.930 136.125 37.335 139.455 ;
        RECT 41.580 133.150 41.950 142.250 ;
        RECT 42.525 134.215 42.815 146.050 ;
        RECT 45.975 144.490 46.385 147.585 ;
        RECT 50.430 143.945 50.740 146.460 ;
        RECT 46.340 136.180 46.780 139.455 ;
        RECT 48.720 138.195 49.245 142.135 ;
        RECT 47.880 134.090 48.205 136.855 ;
        RECT 50.395 136.185 50.810 138.575 ;
        RECT 51.425 134.745 51.740 145.430 ;
        RECT 52.755 139.135 53.240 142.145 ;
        RECT 52.125 133.355 52.460 134.705 ;
        RECT -8.160 117.530 -7.805 131.320 ;
        RECT 55.185 130.690 55.635 140.955 ;
        RECT -6.535 118.385 -6.175 129.720 ;
        RECT 56.350 129.150 56.835 138.035 ;
        RECT 62.655 128.775 63.060 140.305 ;
        RECT 64.730 130.675 65.120 141.775 ;
        RECT 68.500 134.225 68.855 145.310 ;
        RECT 72.245 143.950 72.535 146.010 ;
        RECT 75.015 144.550 75.515 147.600 ;
        RECT 79.985 144.460 80.395 147.555 ;
        RECT 79.025 142.800 79.335 142.830 ;
        RECT 69.825 139.080 70.295 142.070 ;
        RECT 72.175 136.095 72.490 138.465 ;
        RECT 73.795 138.140 74.215 142.105 ;
        RECT 70.460 133.385 70.840 134.760 ;
        RECT 72.900 132.355 73.245 134.815 ;
        RECT 74.535 134.035 74.860 136.800 ;
        RECT 75.520 136.070 75.925 139.400 ;
        RECT 79.025 136.700 79.340 142.800 ;
        RECT 80.170 133.095 80.540 142.195 ;
        RECT 81.115 134.160 81.405 145.995 ;
        RECT 84.565 144.435 84.975 147.530 ;
        RECT 89.020 143.890 89.330 146.405 ;
        RECT 93.270 145.590 93.650 145.970 ;
        RECT 95.400 145.590 95.780 145.970 ;
        RECT 82.010 136.655 82.340 142.850 ;
        RECT 84.915 136.125 85.370 139.400 ;
        RECT 87.275 138.140 87.820 142.080 ;
        RECT 91.330 139.080 91.765 142.090 ;
        RECT 86.470 134.035 86.795 136.800 ;
        RECT 88.985 136.130 89.400 138.520 ;
        RECT 92.525 134.705 92.855 145.400 ;
        RECT 93.960 139.040 94.345 144.825 ;
        RECT 90.715 133.300 91.050 134.650 ;
        RECT 94.320 134.285 94.745 138.560 ;
        RECT 96.020 136.050 96.320 143.090 ;
        RECT 97.140 135.445 97.440 142.375 ;
        RECT 98.450 136.045 98.750 142.395 ;
        RECT 92.980 133.375 93.360 133.755 ;
        RECT 95.175 133.360 95.555 133.740 ;
        RECT 99.045 133.300 99.335 143.080 ;
        RECT 99.765 136.075 100.060 142.900 ;
        RECT 100.895 135.535 101.195 142.345 ;
        RECT 101.685 136.130 101.995 146.170 ;
        RECT 110.875 144.415 111.255 144.795 ;
        RECT 102.480 136.060 102.780 142.890 ;
        RECT 103.605 135.445 103.905 142.385 ;
        RECT 105.055 135.320 105.335 138.355 ;
        RECT 105.815 136.020 106.095 142.380 ;
        RECT 106.665 136.020 106.965 142.840 ;
        RECT 107.805 135.275 108.105 142.430 ;
        RECT 108.450 139.465 108.830 139.845 ;
        RECT 108.450 137.410 108.830 137.790 ;
        RECT 110.300 137.290 110.615 141.615 ;
        RECT 110.910 139.365 111.190 140.895 ;
        RECT 111.480 136.050 111.780 143.090 ;
        RECT 113.255 136.805 113.555 140.865 ;
        RECT 110.775 134.240 111.155 134.620 ;
        RECT 114.505 133.835 114.795 143.080 ;
        RECT 116.355 135.535 116.655 142.345 ;
        RECT 117.145 136.130 117.455 144.865 ;
        RECT 117.940 136.060 118.240 142.890 ;
        RECT 119.745 136.790 120.025 140.880 ;
        RECT 120.515 135.320 120.795 138.355 ;
        RECT 123.265 135.275 123.565 142.430 ;
        RECT -1.050 115.810 -0.750 122.740 ;
        RECT 0.260 116.410 0.560 122.760 ;
        RECT 1.575 116.440 1.870 123.265 ;
        RECT 5.415 115.810 5.715 122.750 ;
        RECT 7.625 116.385 7.930 122.745 ;
        RECT 8.475 116.385 8.775 123.205 ;
        RECT 10.285 119.830 10.665 120.210 ;
        RECT 12.070 118.410 12.390 120.540 ;
        RECT 10.500 115.120 10.880 118.140 ;
        RECT 12.680 117.570 12.960 119.975 ;
        RECT 13.290 116.415 13.590 123.455 ;
        RECT 14.410 115.810 14.710 122.740 ;
        RECT 15.720 116.410 16.020 122.760 ;
        RECT 16.315 118.285 16.640 123.445 ;
        RECT 17.035 116.440 17.330 123.265 ;
        RECT 18.165 115.900 18.465 122.710 ;
        RECT 18.955 116.495 19.265 122.685 ;
        RECT 19.750 116.425 20.050 123.255 ;
        RECT 20.875 115.810 21.175 122.750 ;
        RECT 22.325 115.685 22.605 118.720 ;
        RECT 23.085 116.385 23.405 122.745 ;
        RECT 23.935 116.385 24.235 123.205 ;
        RECT 25.075 115.640 25.375 122.795 ;
        RECT 25.710 117.785 26.090 118.165 ;
        RECT 26.415 113.670 26.775 120.230 ;
        RECT 27.555 118.420 27.880 120.285 ;
        RECT 28.220 115.075 28.680 119.760 ;
        RECT 29.005 117.620 29.455 126.440 ;
        RECT 31.190 119.445 31.620 122.435 ;
        RECT 28.935 113.730 29.315 114.110 ;
        RECT 31.825 113.750 32.205 115.125 ;
        RECT 32.595 114.570 32.910 125.620 ;
        RECT 33.610 124.315 33.900 126.375 ;
        RECT 36.395 124.915 36.870 127.965 ;
        RECT 41.350 124.825 41.760 127.920 ;
        RECT 33.530 116.460 33.855 118.830 ;
        RECT 35.180 118.505 35.580 122.470 ;
        RECT 34.265 112.720 34.610 115.180 ;
        RECT 35.900 114.400 36.225 117.165 ;
        RECT 36.885 116.435 37.290 119.765 ;
        RECT 41.535 113.460 41.905 122.560 ;
        RECT 42.480 114.525 42.770 126.360 ;
        RECT 45.930 124.800 46.340 127.895 ;
        RECT 50.385 124.255 50.695 126.770 ;
        RECT 46.295 116.490 46.735 119.765 ;
        RECT 48.675 118.505 49.200 122.445 ;
        RECT 47.835 114.400 48.160 117.165 ;
        RECT 50.350 116.495 50.765 118.885 ;
        RECT 51.380 115.055 51.695 125.740 ;
        RECT 52.710 119.445 53.195 122.455 ;
        RECT 52.080 113.665 52.415 115.015 ;
        RECT -8.160 97.765 -7.805 111.820 ;
        RECT 55.185 111.190 55.635 121.305 ;
        RECT -6.535 98.570 -6.175 110.220 ;
        RECT 56.350 109.650 56.835 118.405 ;
        RECT 62.955 109.025 63.360 120.555 ;
        RECT 65.030 110.925 65.420 122.025 ;
        RECT 68.300 114.500 68.655 125.585 ;
        RECT 72.045 124.225 72.335 126.285 ;
        RECT 74.815 124.825 75.315 127.875 ;
        RECT 79.785 124.735 80.195 127.830 ;
        RECT 78.825 123.075 79.135 123.105 ;
        RECT 69.625 119.355 70.095 122.345 ;
        RECT 71.975 116.370 72.290 118.740 ;
        RECT 73.595 118.415 74.015 122.380 ;
        RECT 70.260 113.660 70.640 115.035 ;
        RECT 72.700 112.630 73.045 115.090 ;
        RECT 74.335 114.310 74.660 117.075 ;
        RECT 75.320 116.345 75.725 119.675 ;
        RECT 78.825 116.975 79.140 123.075 ;
        RECT 79.970 113.370 80.340 122.470 ;
        RECT 80.915 114.435 81.205 126.270 ;
        RECT 84.365 124.710 84.775 127.805 ;
        RECT 88.820 124.165 89.130 126.680 ;
        RECT 93.070 125.865 93.450 126.245 ;
        RECT 95.200 125.865 95.580 126.245 ;
        RECT 81.810 116.930 82.140 123.125 ;
        RECT 84.715 116.400 85.170 119.675 ;
        RECT 87.075 118.415 87.620 122.355 ;
        RECT 91.130 119.355 91.565 122.365 ;
        RECT 86.270 114.310 86.595 117.075 ;
        RECT 88.785 116.405 89.200 118.795 ;
        RECT 92.325 114.980 92.655 125.675 ;
        RECT 93.760 119.315 94.145 125.100 ;
        RECT 90.515 113.575 90.850 114.925 ;
        RECT 94.120 114.560 94.545 118.835 ;
        RECT 95.820 116.325 96.120 123.365 ;
        RECT 96.940 115.720 97.240 122.650 ;
        RECT 98.250 116.320 98.550 122.670 ;
        RECT 92.780 113.650 93.160 114.030 ;
        RECT 94.975 113.635 95.355 114.015 ;
        RECT 98.845 113.575 99.135 123.355 ;
        RECT 99.565 116.350 99.860 123.175 ;
        RECT 100.695 115.810 100.995 122.620 ;
        RECT 101.485 116.405 101.795 126.445 ;
        RECT 110.675 124.690 111.055 125.070 ;
        RECT 102.280 116.335 102.580 123.165 ;
        RECT 103.405 115.720 103.705 122.660 ;
        RECT 104.855 115.595 105.135 118.630 ;
        RECT 105.615 116.295 105.895 122.655 ;
        RECT 106.465 116.295 106.765 123.115 ;
        RECT 107.605 115.550 107.905 122.705 ;
        RECT 108.250 119.740 108.630 120.120 ;
        RECT 108.250 117.685 108.630 118.065 ;
        RECT 110.100 117.565 110.415 121.890 ;
        RECT 110.710 119.640 110.990 121.170 ;
        RECT 111.280 116.325 111.580 123.365 ;
        RECT 113.055 117.080 113.355 121.140 ;
        RECT 110.575 114.515 110.955 114.895 ;
        RECT 114.305 114.110 114.595 123.355 ;
        RECT 116.155 115.810 116.455 122.620 ;
        RECT 116.945 116.405 117.255 125.140 ;
        RECT 117.740 116.335 118.040 123.165 ;
        RECT 119.545 117.065 119.825 121.155 ;
        RECT 120.315 115.595 120.595 118.630 ;
        RECT 123.065 115.550 123.365 122.705 ;
        RECT 125.105 121.445 125.480 129.645 ;
        RECT 126.850 120.640 127.150 131.635 ;
        RECT -0.860 96.100 -0.560 103.030 ;
        RECT 0.450 96.700 0.750 103.050 ;
        RECT 1.765 96.730 2.060 103.555 ;
        RECT 5.605 96.100 5.905 103.040 ;
        RECT 7.815 96.675 8.120 103.035 ;
        RECT 8.665 96.675 8.965 103.495 ;
        RECT 10.475 100.120 10.855 100.500 ;
        RECT 12.260 98.700 12.580 100.830 ;
        RECT 10.690 95.410 11.070 98.430 ;
        RECT 12.870 97.860 13.150 100.265 ;
        RECT 13.480 96.705 13.780 103.745 ;
        RECT 14.600 96.100 14.900 103.030 ;
        RECT 15.910 96.700 16.210 103.050 ;
        RECT 16.505 98.575 16.830 103.735 ;
        RECT 17.225 96.730 17.520 103.555 ;
        RECT 18.355 96.190 18.655 103.000 ;
        RECT 19.145 96.785 19.455 102.975 ;
        RECT 19.940 96.715 20.240 103.545 ;
        RECT 21.065 96.100 21.365 103.040 ;
        RECT 22.515 95.975 22.795 99.010 ;
        RECT 23.275 96.675 23.595 103.035 ;
        RECT 24.125 96.675 24.425 103.495 ;
        RECT 25.265 95.930 25.565 103.085 ;
        RECT 25.900 98.075 26.280 98.455 ;
        RECT 26.605 93.960 26.965 100.520 ;
        RECT 27.745 98.710 28.070 100.575 ;
        RECT 28.410 95.365 28.870 100.050 ;
        RECT 29.195 97.910 29.645 106.730 ;
        RECT 31.380 99.735 31.810 102.725 ;
        RECT 29.125 94.020 29.505 94.400 ;
        RECT 32.015 94.040 32.395 95.415 ;
        RECT 32.785 94.860 33.100 105.910 ;
        RECT 33.800 104.605 34.090 106.665 ;
        RECT 36.585 105.205 37.060 108.255 ;
        RECT 41.540 105.115 41.950 108.210 ;
        RECT 33.720 96.750 34.045 99.120 ;
        RECT 35.370 98.795 35.770 102.760 ;
        RECT 34.455 93.010 34.800 95.470 ;
        RECT 36.090 94.690 36.415 97.455 ;
        RECT 37.075 96.725 37.480 100.055 ;
        RECT 41.725 93.750 42.095 102.850 ;
        RECT 42.670 94.815 42.960 106.650 ;
        RECT 46.120 105.090 46.530 108.185 ;
        RECT 50.575 104.545 50.885 107.060 ;
        RECT 46.485 96.780 46.925 100.055 ;
        RECT 48.865 98.795 49.390 102.735 ;
        RECT 48.025 94.690 48.350 97.455 ;
        RECT 50.540 96.785 50.955 99.175 ;
        RECT 51.570 95.345 51.885 106.030 ;
        RECT 52.900 99.735 53.385 102.745 ;
        RECT 52.270 93.955 52.605 95.305 ;
        RECT -7.950 77.990 -7.595 91.780 ;
        RECT 55.395 91.150 55.845 101.650 ;
        RECT -6.325 78.845 -5.965 90.180 ;
        RECT 56.560 89.610 57.045 98.850 ;
        RECT 62.975 89.365 63.380 100.895 ;
        RECT 65.050 91.265 65.440 102.365 ;
        RECT 68.455 94.855 68.810 105.940 ;
        RECT 72.200 104.580 72.490 106.640 ;
        RECT 74.970 105.180 75.470 108.230 ;
        RECT 79.940 105.090 80.350 108.185 ;
        RECT 78.980 103.430 79.290 103.460 ;
        RECT 69.780 99.710 70.250 102.700 ;
        RECT 72.130 96.725 72.445 99.095 ;
        RECT 73.750 98.770 74.170 102.735 ;
        RECT 70.415 94.015 70.795 95.390 ;
        RECT 72.855 92.985 73.200 95.445 ;
        RECT 74.490 94.665 74.815 97.430 ;
        RECT 75.475 96.700 75.880 100.030 ;
        RECT 78.980 97.330 79.295 103.430 ;
        RECT 80.125 93.725 80.495 102.825 ;
        RECT 81.070 94.790 81.360 106.625 ;
        RECT 84.520 105.065 84.930 108.160 ;
        RECT 88.975 104.520 89.285 107.035 ;
        RECT 93.225 106.220 93.605 106.600 ;
        RECT 95.355 106.220 95.735 106.600 ;
        RECT 81.965 97.285 82.295 103.480 ;
        RECT 84.870 96.755 85.325 100.030 ;
        RECT 87.230 98.770 87.775 102.710 ;
        RECT 91.285 99.710 91.720 102.720 ;
        RECT 86.425 94.665 86.750 97.430 ;
        RECT 88.940 96.760 89.355 99.150 ;
        RECT 92.480 95.335 92.810 106.030 ;
        RECT 93.915 99.670 94.300 105.455 ;
        RECT 90.670 93.930 91.005 95.280 ;
        RECT 94.275 94.915 94.700 99.190 ;
        RECT 95.975 96.680 96.275 103.720 ;
        RECT 97.095 96.075 97.395 103.005 ;
        RECT 98.405 96.675 98.705 103.025 ;
        RECT 92.935 94.005 93.315 94.385 ;
        RECT 95.130 93.990 95.510 94.370 ;
        RECT 99.000 93.930 99.290 103.710 ;
        RECT 99.720 96.705 100.015 103.530 ;
        RECT 100.850 96.165 101.150 102.975 ;
        RECT 101.640 96.760 101.950 106.800 ;
        RECT 110.830 105.045 111.210 105.425 ;
        RECT 102.435 96.690 102.735 103.520 ;
        RECT 103.560 96.075 103.860 103.015 ;
        RECT 105.010 95.950 105.290 98.985 ;
        RECT 105.770 96.650 106.050 103.010 ;
        RECT 106.620 96.650 106.920 103.470 ;
        RECT 107.760 95.905 108.060 103.060 ;
        RECT 108.405 100.095 108.785 100.475 ;
        RECT 108.405 98.040 108.785 98.420 ;
        RECT 110.255 97.920 110.570 102.245 ;
        RECT 110.865 99.995 111.145 101.525 ;
        RECT 111.435 96.680 111.735 103.720 ;
        RECT 113.210 97.435 113.510 101.495 ;
        RECT 110.730 94.870 111.110 95.250 ;
        RECT 114.460 94.465 114.750 103.710 ;
        RECT 116.310 96.165 116.610 102.975 ;
        RECT 117.100 96.760 117.410 105.495 ;
        RECT 117.895 96.690 118.195 103.520 ;
        RECT 119.700 97.420 119.980 101.510 ;
        RECT 120.470 95.950 120.750 98.985 ;
        RECT 123.220 95.905 123.520 103.060 ;
        RECT 125.405 101.695 125.780 109.895 ;
        RECT 127.150 100.890 127.450 111.885 ;
        RECT -1.055 76.260 -0.755 83.190 ;
        RECT 0.255 76.860 0.555 83.210 ;
        RECT 1.570 76.890 1.865 83.715 ;
        RECT 5.410 76.260 5.710 83.200 ;
        RECT 7.620 76.835 7.925 83.195 ;
        RECT 8.470 76.835 8.770 83.655 ;
        RECT 10.280 80.280 10.660 80.660 ;
        RECT 12.065 78.860 12.385 80.990 ;
        RECT 10.495 75.570 10.875 78.590 ;
        RECT 12.675 78.020 12.955 80.425 ;
        RECT 13.285 76.865 13.585 83.905 ;
        RECT 14.405 76.260 14.705 83.190 ;
        RECT 15.715 76.860 16.015 83.210 ;
        RECT 16.310 78.735 16.635 83.895 ;
        RECT 17.030 76.890 17.325 83.715 ;
        RECT 18.160 76.350 18.460 83.160 ;
        RECT 18.950 76.945 19.260 83.135 ;
        RECT 19.745 76.875 20.045 83.705 ;
        RECT 20.870 76.260 21.170 83.200 ;
        RECT 22.320 76.135 22.600 79.170 ;
        RECT 23.080 76.835 23.400 83.195 ;
        RECT 23.930 76.835 24.230 83.655 ;
        RECT 25.070 76.090 25.370 83.245 ;
        RECT 25.705 78.235 26.085 78.615 ;
        RECT 26.410 74.120 26.770 80.680 ;
        RECT 27.550 78.870 27.875 80.735 ;
        RECT 28.215 75.525 28.675 80.210 ;
        RECT 29.000 78.070 29.450 86.890 ;
        RECT 31.185 79.895 31.615 82.885 ;
        RECT 28.930 74.180 29.310 74.560 ;
        RECT 31.820 74.200 32.200 75.575 ;
        RECT 32.590 75.020 32.905 86.070 ;
        RECT 33.605 84.765 33.895 86.825 ;
        RECT 36.390 85.365 36.865 88.415 ;
        RECT 41.345 85.275 41.755 88.370 ;
        RECT 33.525 76.910 33.850 79.280 ;
        RECT 35.175 78.955 35.575 82.920 ;
        RECT 34.260 73.170 34.605 75.630 ;
        RECT 35.895 74.850 36.220 77.615 ;
        RECT 36.880 76.885 37.285 80.215 ;
        RECT 41.530 73.910 41.900 83.010 ;
        RECT 42.475 74.975 42.765 86.810 ;
        RECT 45.925 85.250 46.335 88.345 ;
        RECT 50.380 84.705 50.690 87.220 ;
        RECT 46.290 76.940 46.730 80.215 ;
        RECT 48.670 78.955 49.195 82.895 ;
        RECT 47.830 74.850 48.155 77.615 ;
        RECT 50.345 76.945 50.760 79.335 ;
        RECT 51.375 75.505 51.690 86.190 ;
        RECT 52.705 79.895 53.190 82.905 ;
        RECT 52.075 74.115 52.410 75.465 ;
        RECT -7.995 58.200 -7.640 71.990 ;
        RECT 55.350 71.360 55.800 81.850 ;
        RECT -6.370 59.105 -6.010 70.390 ;
        RECT 56.515 69.820 57.000 78.980 ;
        RECT 62.975 69.630 63.380 81.160 ;
        RECT 65.050 71.530 65.440 82.630 ;
        RECT 68.455 75.060 68.810 86.145 ;
        RECT 72.200 84.785 72.490 86.845 ;
        RECT 74.970 85.385 75.470 88.435 ;
        RECT 79.940 85.295 80.350 88.390 ;
        RECT 78.980 83.635 79.290 83.665 ;
        RECT 69.780 79.915 70.250 82.905 ;
        RECT 72.130 76.930 72.445 79.300 ;
        RECT 73.750 78.975 74.170 82.940 ;
        RECT 70.415 74.220 70.795 75.595 ;
        RECT 72.855 73.190 73.200 75.650 ;
        RECT 74.490 74.870 74.815 77.635 ;
        RECT 75.475 76.905 75.880 80.235 ;
        RECT 78.980 77.535 79.295 83.635 ;
        RECT 80.125 73.930 80.495 83.030 ;
        RECT 81.070 74.995 81.360 86.830 ;
        RECT 84.520 85.270 84.930 88.365 ;
        RECT 88.975 84.725 89.285 87.240 ;
        RECT 93.225 86.425 93.605 86.805 ;
        RECT 95.355 86.425 95.735 86.805 ;
        RECT 81.965 77.490 82.295 83.685 ;
        RECT 84.870 76.960 85.325 80.235 ;
        RECT 87.230 78.975 87.775 82.915 ;
        RECT 91.285 79.915 91.720 82.925 ;
        RECT 86.425 74.870 86.750 77.635 ;
        RECT 88.940 76.965 89.355 79.355 ;
        RECT 92.480 75.540 92.810 86.235 ;
        RECT 93.915 79.875 94.300 85.660 ;
        RECT 90.670 74.135 91.005 75.485 ;
        RECT 94.275 75.120 94.700 79.395 ;
        RECT 95.975 76.885 96.275 83.925 ;
        RECT 97.095 76.280 97.395 83.210 ;
        RECT 98.405 76.880 98.705 83.230 ;
        RECT 92.935 74.210 93.315 74.590 ;
        RECT 95.130 74.195 95.510 74.575 ;
        RECT 99.000 74.135 99.290 83.915 ;
        RECT 99.720 76.910 100.015 83.735 ;
        RECT 100.850 76.370 101.150 83.180 ;
        RECT 101.640 76.965 101.950 87.005 ;
        RECT 110.830 85.250 111.210 85.630 ;
        RECT 102.435 76.895 102.735 83.725 ;
        RECT 103.560 76.280 103.860 83.220 ;
        RECT 105.010 76.155 105.290 79.190 ;
        RECT 105.770 76.855 106.050 83.215 ;
        RECT 106.620 76.855 106.920 83.675 ;
        RECT 107.760 76.110 108.060 83.265 ;
        RECT 108.405 80.300 108.785 80.680 ;
        RECT 108.405 78.245 108.785 78.625 ;
        RECT 110.255 78.125 110.570 82.450 ;
        RECT 110.865 80.200 111.145 81.730 ;
        RECT 111.435 76.885 111.735 83.925 ;
        RECT 113.210 77.640 113.510 81.700 ;
        RECT 110.730 75.075 111.110 75.455 ;
        RECT 114.460 74.670 114.750 83.915 ;
        RECT 116.310 76.370 116.610 83.180 ;
        RECT 117.100 76.965 117.410 85.700 ;
        RECT 117.895 76.895 118.195 83.725 ;
        RECT 119.700 77.625 119.980 81.715 ;
        RECT 120.470 76.155 120.750 79.190 ;
        RECT 123.220 76.110 123.520 83.265 ;
        RECT 125.425 82.035 125.800 90.235 ;
        RECT 127.170 81.230 127.470 92.225 ;
        RECT -1.185 56.550 -0.885 63.480 ;
        RECT 0.125 57.150 0.425 63.500 ;
        RECT 1.440 57.180 1.735 64.005 ;
        RECT 5.280 56.550 5.580 63.490 ;
        RECT 7.490 57.125 7.795 63.485 ;
        RECT 8.340 57.125 8.640 63.945 ;
        RECT 10.150 60.570 10.530 60.950 ;
        RECT 11.935 59.150 12.255 61.280 ;
        RECT 10.365 55.860 10.745 58.880 ;
        RECT 12.545 58.310 12.825 60.715 ;
        RECT 13.155 57.155 13.455 64.195 ;
        RECT 14.275 56.550 14.575 63.480 ;
        RECT 15.585 57.150 15.885 63.500 ;
        RECT 16.180 59.025 16.505 64.185 ;
        RECT 16.900 57.180 17.195 64.005 ;
        RECT 18.030 56.640 18.330 63.450 ;
        RECT 18.820 57.235 19.130 63.425 ;
        RECT 19.615 57.165 19.915 63.995 ;
        RECT 20.740 56.550 21.040 63.490 ;
        RECT 22.190 56.425 22.470 59.460 ;
        RECT 22.950 57.125 23.270 63.485 ;
        RECT 23.800 57.125 24.100 63.945 ;
        RECT 24.940 56.380 25.240 63.535 ;
        RECT 25.575 58.525 25.955 58.905 ;
        RECT 26.280 54.410 26.640 60.970 ;
        RECT 27.420 59.160 27.745 61.025 ;
        RECT 28.085 55.815 28.545 60.500 ;
        RECT 28.870 58.360 29.320 67.180 ;
        RECT 31.055 60.185 31.485 63.175 ;
        RECT 28.800 54.470 29.180 54.850 ;
        RECT 31.690 54.490 32.070 55.865 ;
        RECT 32.460 55.310 32.775 66.360 ;
        RECT 33.475 65.055 33.765 67.115 ;
        RECT 36.260 65.655 36.735 68.705 ;
        RECT 41.215 65.565 41.625 68.660 ;
        RECT 33.395 57.200 33.720 59.570 ;
        RECT 35.045 59.245 35.445 63.210 ;
        RECT 34.130 53.460 34.475 55.920 ;
        RECT 35.765 55.140 36.090 57.905 ;
        RECT 36.750 57.175 37.155 60.505 ;
        RECT 41.400 54.200 41.770 63.300 ;
        RECT 42.345 55.265 42.635 67.100 ;
        RECT 45.795 65.540 46.205 68.635 ;
        RECT 50.250 64.995 50.560 67.510 ;
        RECT 46.160 57.230 46.600 60.505 ;
        RECT 48.540 59.245 49.065 63.185 ;
        RECT 47.700 55.140 48.025 57.905 ;
        RECT 50.215 57.235 50.630 59.625 ;
        RECT 51.245 55.795 51.560 66.480 ;
        RECT 52.575 60.185 53.060 63.195 ;
        RECT 51.945 54.405 52.280 55.755 ;
        RECT -8.300 38.440 -7.945 52.360 ;
        RECT 55.045 51.730 55.495 61.995 ;
        RECT -6.675 39.345 -6.315 50.760 ;
        RECT 56.210 50.190 56.695 59.075 ;
        RECT 62.875 49.925 63.280 61.455 ;
        RECT 64.950 51.825 65.340 62.925 ;
        RECT 68.375 55.305 68.730 66.390 ;
        RECT 72.120 65.030 72.410 67.090 ;
        RECT 74.890 65.630 75.390 68.680 ;
        RECT 79.860 65.540 80.270 68.635 ;
        RECT 78.900 63.880 79.210 63.910 ;
        RECT 69.700 60.160 70.170 63.150 ;
        RECT 72.050 57.175 72.365 59.545 ;
        RECT 73.670 59.220 74.090 63.185 ;
        RECT 70.335 54.465 70.715 55.840 ;
        RECT 72.775 53.435 73.120 55.895 ;
        RECT 74.410 55.115 74.735 57.880 ;
        RECT 75.395 57.150 75.800 60.480 ;
        RECT 78.900 57.780 79.215 63.880 ;
        RECT 80.045 54.175 80.415 63.275 ;
        RECT 80.990 55.240 81.280 67.075 ;
        RECT 84.440 65.515 84.850 68.610 ;
        RECT 88.895 64.970 89.205 67.485 ;
        RECT 93.145 66.670 93.525 67.050 ;
        RECT 95.275 66.670 95.655 67.050 ;
        RECT 81.885 57.735 82.215 63.930 ;
        RECT 84.790 57.205 85.245 60.480 ;
        RECT 87.150 59.220 87.695 63.160 ;
        RECT 91.205 60.160 91.640 63.170 ;
        RECT 86.345 55.115 86.670 57.880 ;
        RECT 88.860 57.210 89.275 59.600 ;
        RECT 92.400 55.785 92.730 66.480 ;
        RECT 93.835 60.120 94.220 65.905 ;
        RECT 90.590 54.380 90.925 55.730 ;
        RECT 94.195 55.365 94.620 59.640 ;
        RECT 95.895 57.130 96.195 64.170 ;
        RECT 97.015 56.525 97.315 63.455 ;
        RECT 98.325 57.125 98.625 63.475 ;
        RECT 92.855 54.455 93.235 54.835 ;
        RECT 95.050 54.440 95.430 54.820 ;
        RECT 98.920 54.380 99.210 64.160 ;
        RECT 99.640 57.155 99.935 63.980 ;
        RECT 100.770 56.615 101.070 63.425 ;
        RECT 101.560 57.210 101.870 67.250 ;
        RECT 110.750 65.495 111.130 65.875 ;
        RECT 102.355 57.140 102.655 63.970 ;
        RECT 103.480 56.525 103.780 63.465 ;
        RECT 104.930 56.400 105.210 59.435 ;
        RECT 105.690 57.100 105.970 63.460 ;
        RECT 106.540 57.100 106.840 63.920 ;
        RECT 107.680 56.355 107.980 63.510 ;
        RECT 108.325 60.545 108.705 60.925 ;
        RECT 108.325 58.490 108.705 58.870 ;
        RECT 110.175 58.370 110.490 62.695 ;
        RECT 110.785 60.445 111.065 61.975 ;
        RECT 111.355 57.130 111.655 64.170 ;
        RECT 113.130 57.885 113.430 61.945 ;
        RECT 110.650 55.320 111.030 55.700 ;
        RECT 114.380 54.915 114.670 64.160 ;
        RECT 116.230 56.615 116.530 63.425 ;
        RECT 117.020 57.210 117.330 65.945 ;
        RECT 117.815 57.140 118.115 63.970 ;
        RECT 119.620 57.870 119.900 61.960 ;
        RECT 120.390 56.400 120.670 59.435 ;
        RECT 123.140 56.355 123.440 63.510 ;
        RECT 125.425 62.215 125.800 70.500 ;
        RECT 127.170 61.495 127.470 72.490 ;
        RECT -1.055 36.790 -0.755 43.720 ;
        RECT 0.255 37.390 0.555 43.740 ;
        RECT 1.570 37.420 1.865 44.245 ;
        RECT 5.410 36.790 5.710 43.730 ;
        RECT 7.620 37.365 7.925 43.725 ;
        RECT 8.470 37.365 8.770 44.185 ;
        RECT 10.280 40.810 10.660 41.190 ;
        RECT 12.065 39.390 12.385 41.520 ;
        RECT 10.495 36.100 10.875 39.120 ;
        RECT 12.675 38.550 12.955 40.955 ;
        RECT 13.285 37.395 13.585 44.435 ;
        RECT 14.405 36.790 14.705 43.720 ;
        RECT 15.715 37.390 16.015 43.740 ;
        RECT 16.310 39.265 16.635 44.425 ;
        RECT 17.030 37.420 17.325 44.245 ;
        RECT 18.160 36.880 18.460 43.690 ;
        RECT 18.950 37.475 19.260 43.665 ;
        RECT 19.745 37.405 20.045 44.235 ;
        RECT 20.870 36.790 21.170 43.730 ;
        RECT 22.320 36.665 22.600 39.700 ;
        RECT 23.080 37.365 23.400 43.725 ;
        RECT 23.930 37.365 24.230 44.185 ;
        RECT 25.070 36.620 25.370 43.775 ;
        RECT 25.705 38.765 26.085 39.145 ;
        RECT 26.410 34.650 26.770 41.210 ;
        RECT 27.550 39.400 27.875 41.265 ;
        RECT 28.215 36.055 28.675 40.740 ;
        RECT 29.000 38.600 29.450 47.420 ;
        RECT 31.185 40.425 31.615 43.415 ;
        RECT 28.930 34.710 29.310 35.090 ;
        RECT 31.820 34.730 32.200 36.105 ;
        RECT 32.590 35.550 32.905 46.600 ;
        RECT 33.605 45.295 33.895 47.355 ;
        RECT 36.390 45.895 36.865 48.945 ;
        RECT 41.345 45.805 41.755 48.900 ;
        RECT 33.525 37.440 33.850 39.810 ;
        RECT 35.175 39.485 35.575 43.450 ;
        RECT 34.260 33.700 34.605 36.160 ;
        RECT 35.895 35.380 36.220 38.145 ;
        RECT 36.880 37.415 37.285 40.745 ;
        RECT 41.530 34.440 41.900 43.540 ;
        RECT 42.475 35.505 42.765 47.340 ;
        RECT 45.925 45.780 46.335 48.875 ;
        RECT 50.380 45.235 50.690 47.750 ;
        RECT 46.290 37.470 46.730 40.745 ;
        RECT 48.670 39.485 49.195 43.425 ;
        RECT 47.830 35.380 48.155 38.145 ;
        RECT 50.345 37.475 50.760 39.865 ;
        RECT 51.375 36.035 51.690 46.720 ;
        RECT 52.705 40.425 53.190 43.435 ;
        RECT 52.075 34.645 52.410 35.995 ;
        RECT -8.205 18.675 -7.850 32.585 ;
        RECT 55.140 31.955 55.590 42.220 ;
        RECT -6.580 19.595 -6.220 30.985 ;
        RECT 56.305 30.415 56.790 39.300 ;
        RECT 63.135 29.770 63.540 41.650 ;
        RECT 65.210 31.670 65.600 43.250 ;
        RECT 68.480 35.590 68.835 46.675 ;
        RECT 72.225 45.315 72.515 47.375 ;
        RECT 74.995 45.915 75.495 48.965 ;
        RECT 79.965 45.825 80.375 48.920 ;
        RECT 79.005 44.165 79.315 44.195 ;
        RECT 69.805 40.445 70.275 43.435 ;
        RECT 72.155 37.460 72.470 39.830 ;
        RECT 73.775 39.505 74.195 43.470 ;
        RECT 70.440 34.750 70.820 36.125 ;
        RECT 72.880 33.720 73.225 36.180 ;
        RECT 74.515 35.400 74.840 38.165 ;
        RECT 75.500 37.435 75.905 40.765 ;
        RECT 79.005 38.065 79.320 44.165 ;
        RECT 80.150 34.460 80.520 43.560 ;
        RECT 81.095 35.525 81.385 47.360 ;
        RECT 84.545 45.800 84.955 48.895 ;
        RECT 89.000 45.255 89.310 47.770 ;
        RECT 93.250 46.955 93.630 47.335 ;
        RECT 95.380 46.955 95.760 47.335 ;
        RECT 81.990 38.020 82.320 44.215 ;
        RECT 84.895 37.490 85.350 40.765 ;
        RECT 87.255 39.505 87.800 43.445 ;
        RECT 91.310 40.445 91.745 43.455 ;
        RECT 86.450 35.400 86.775 38.165 ;
        RECT 88.965 37.495 89.380 39.885 ;
        RECT 92.505 36.070 92.835 46.765 ;
        RECT 93.940 40.405 94.325 46.190 ;
        RECT 90.695 34.665 91.030 36.015 ;
        RECT 94.300 35.650 94.725 39.925 ;
        RECT 96.000 37.415 96.300 44.455 ;
        RECT 97.120 36.810 97.420 43.740 ;
        RECT 98.430 37.410 98.730 43.760 ;
        RECT 92.960 34.740 93.340 35.120 ;
        RECT 95.155 34.725 95.535 35.105 ;
        RECT 99.025 34.665 99.315 44.445 ;
        RECT 99.745 37.440 100.040 44.265 ;
        RECT 100.875 36.900 101.175 43.710 ;
        RECT 101.665 37.495 101.975 47.535 ;
        RECT 110.855 45.780 111.235 46.160 ;
        RECT 102.460 37.425 102.760 44.255 ;
        RECT 103.585 36.810 103.885 43.750 ;
        RECT 105.035 36.685 105.315 39.720 ;
        RECT 105.795 37.385 106.075 43.745 ;
        RECT 106.645 37.385 106.945 44.205 ;
        RECT 107.785 36.640 108.085 43.795 ;
        RECT 108.430 40.830 108.810 41.210 ;
        RECT 108.430 38.775 108.810 39.155 ;
        RECT 110.280 38.655 110.595 42.980 ;
        RECT 110.890 40.730 111.170 42.260 ;
        RECT 111.460 37.415 111.760 44.455 ;
        RECT 113.235 38.170 113.535 42.230 ;
        RECT 110.755 35.605 111.135 35.985 ;
        RECT 114.485 35.200 114.775 44.445 ;
        RECT 116.335 36.900 116.635 43.710 ;
        RECT 117.125 37.495 117.435 46.230 ;
        RECT 117.920 37.425 118.220 44.255 ;
        RECT 119.725 38.155 120.005 42.245 ;
        RECT 120.495 36.685 120.775 39.720 ;
        RECT 123.245 36.640 123.545 43.795 ;
        RECT 125.325 42.515 125.700 50.795 ;
        RECT 127.070 41.675 127.370 52.785 ;
        RECT -1.105 16.980 -0.805 23.910 ;
        RECT 0.205 17.580 0.505 23.930 ;
        RECT 1.520 17.610 1.815 24.435 ;
        RECT 5.360 16.980 5.660 23.920 ;
        RECT 7.570 17.555 7.875 23.915 ;
        RECT 8.420 17.555 8.720 24.375 ;
        RECT 10.230 21.000 10.610 21.380 ;
        RECT 12.015 19.580 12.335 21.710 ;
        RECT 10.445 16.290 10.825 19.310 ;
        RECT 12.625 18.740 12.905 21.145 ;
        RECT 13.235 17.585 13.535 24.625 ;
        RECT 14.355 16.980 14.655 23.910 ;
        RECT 15.665 17.580 15.965 23.930 ;
        RECT 16.260 19.455 16.585 24.615 ;
        RECT 16.980 17.610 17.275 24.435 ;
        RECT 18.110 17.070 18.410 23.880 ;
        RECT 18.900 17.665 19.210 23.855 ;
        RECT 19.695 17.595 19.995 24.425 ;
        RECT 20.820 16.980 21.120 23.920 ;
        RECT 22.270 16.855 22.550 19.890 ;
        RECT 23.030 17.555 23.350 23.915 ;
        RECT 23.880 17.555 24.180 24.375 ;
        RECT 25.020 16.810 25.320 23.965 ;
        RECT 25.655 18.955 26.035 19.335 ;
        RECT 26.360 14.840 26.720 21.400 ;
        RECT 27.500 19.590 27.825 21.455 ;
        RECT 28.165 16.245 28.625 20.930 ;
        RECT 28.950 18.790 29.400 27.610 ;
        RECT 31.135 20.615 31.565 23.605 ;
        RECT 28.880 14.900 29.260 15.280 ;
        RECT 31.770 14.920 32.150 16.295 ;
        RECT 32.540 15.740 32.855 26.790 ;
        RECT 33.555 25.485 33.845 27.545 ;
        RECT 36.340 26.085 36.815 29.135 ;
        RECT 41.295 25.995 41.705 29.090 ;
        RECT 33.475 17.630 33.800 20.000 ;
        RECT 35.125 19.675 35.525 23.640 ;
        RECT 34.210 13.890 34.555 16.350 ;
        RECT 35.845 15.570 36.170 18.335 ;
        RECT 36.830 17.605 37.235 20.935 ;
        RECT 41.480 14.630 41.850 23.730 ;
        RECT 42.425 15.695 42.715 27.530 ;
        RECT 45.875 25.970 46.285 29.065 ;
        RECT 50.330 25.425 50.640 27.940 ;
        RECT 46.240 17.660 46.680 20.935 ;
        RECT 48.620 19.675 49.145 23.615 ;
        RECT 47.780 15.570 48.105 18.335 ;
        RECT 50.295 17.665 50.710 20.055 ;
        RECT 51.325 16.225 51.640 26.910 ;
        RECT 52.655 20.615 53.140 23.625 ;
        RECT 52.025 14.835 52.360 16.185 ;
        RECT -8.205 -1.165 -7.850 12.775 ;
        RECT 55.140 12.145 55.590 22.410 ;
        RECT -6.580 -0.375 -6.220 11.175 ;
        RECT 56.305 10.605 56.790 19.490 ;
        RECT 63.245 9.880 63.650 21.925 ;
        RECT 65.320 11.780 65.710 23.205 ;
        RECT 68.480 15.620 68.835 26.705 ;
        RECT 72.225 25.345 72.515 27.405 ;
        RECT 74.995 25.945 75.495 28.995 ;
        RECT 79.965 25.855 80.375 28.950 ;
        RECT 79.005 24.195 79.315 24.225 ;
        RECT 69.805 20.475 70.275 23.465 ;
        RECT 72.155 17.490 72.470 19.860 ;
        RECT 73.775 19.535 74.195 23.500 ;
        RECT 70.440 14.780 70.820 16.155 ;
        RECT 72.880 13.750 73.225 16.210 ;
        RECT 74.515 15.430 74.840 18.195 ;
        RECT 75.500 17.465 75.905 20.795 ;
        RECT 79.005 18.095 79.320 24.195 ;
        RECT 80.150 14.490 80.520 23.590 ;
        RECT 81.095 15.555 81.385 27.390 ;
        RECT 84.545 25.830 84.955 28.925 ;
        RECT 89.000 25.285 89.310 27.800 ;
        RECT 93.250 26.985 93.630 27.365 ;
        RECT 95.380 26.985 95.760 27.365 ;
        RECT 81.990 18.050 82.320 24.245 ;
        RECT 84.895 17.520 85.350 20.795 ;
        RECT 87.255 19.535 87.800 23.475 ;
        RECT 91.310 20.475 91.745 23.485 ;
        RECT 86.450 15.430 86.775 18.195 ;
        RECT 88.965 17.525 89.380 19.915 ;
        RECT 92.505 16.100 92.835 26.795 ;
        RECT 93.940 20.435 94.325 26.220 ;
        RECT 90.695 14.695 91.030 16.045 ;
        RECT 94.300 15.680 94.725 19.955 ;
        RECT 96.000 17.445 96.300 24.485 ;
        RECT 97.120 16.840 97.420 23.770 ;
        RECT 98.430 17.440 98.730 23.790 ;
        RECT 92.960 14.770 93.340 15.150 ;
        RECT 95.155 14.755 95.535 15.135 ;
        RECT 99.025 14.695 99.315 24.475 ;
        RECT 99.745 17.470 100.040 24.295 ;
        RECT 100.875 16.930 101.175 23.740 ;
        RECT 101.665 17.525 101.975 27.565 ;
        RECT 110.855 25.810 111.235 26.190 ;
        RECT 102.460 17.455 102.760 24.285 ;
        RECT 103.585 16.840 103.885 23.780 ;
        RECT 105.035 16.715 105.315 19.750 ;
        RECT 105.795 17.415 106.075 23.775 ;
        RECT 106.645 17.415 106.945 24.235 ;
        RECT 107.785 16.670 108.085 23.825 ;
        RECT 108.430 20.860 108.810 21.240 ;
        RECT 108.430 18.805 108.810 19.185 ;
        RECT 110.280 18.685 110.595 23.010 ;
        RECT 110.890 20.760 111.170 22.290 ;
        RECT 111.460 17.445 111.760 24.485 ;
        RECT 113.235 18.200 113.535 22.260 ;
        RECT 110.755 15.635 111.135 16.015 ;
        RECT 114.485 15.230 114.775 24.475 ;
        RECT 116.335 16.930 116.635 23.740 ;
        RECT 117.125 17.525 117.435 26.260 ;
        RECT 117.920 17.455 118.220 24.285 ;
        RECT 119.725 18.185 120.005 22.275 ;
        RECT 120.495 16.715 120.775 19.750 ;
        RECT 123.245 16.670 123.545 23.825 ;
        RECT 125.585 22.440 125.960 30.640 ;
        RECT 127.330 21.635 127.630 32.630 ;
        RECT -1.135 -2.815 -0.835 4.115 ;
        RECT 0.175 -2.215 0.475 4.135 ;
        RECT 1.490 -2.185 1.785 4.640 ;
        RECT 5.330 -2.815 5.630 4.125 ;
        RECT 7.540 -2.240 7.845 4.120 ;
        RECT 8.390 -2.240 8.690 4.580 ;
        RECT 10.200 1.205 10.580 1.585 ;
        RECT 11.985 -0.215 12.305 1.915 ;
        RECT 10.415 -3.505 10.795 -0.485 ;
        RECT 12.595 -1.055 12.875 1.350 ;
        RECT 13.205 -2.210 13.505 4.830 ;
        RECT 14.325 -2.815 14.625 4.115 ;
        RECT 15.635 -2.215 15.935 4.135 ;
        RECT 16.230 -0.340 16.555 4.820 ;
        RECT 16.950 -2.185 17.245 4.640 ;
        RECT 18.080 -2.725 18.380 4.085 ;
        RECT 18.870 -2.130 19.180 4.060 ;
        RECT 19.665 -2.200 19.965 4.630 ;
        RECT 20.790 -2.815 21.090 4.125 ;
        RECT 22.240 -2.940 22.520 0.095 ;
        RECT 23.000 -2.240 23.320 4.120 ;
        RECT 23.850 -2.240 24.150 4.580 ;
        RECT 24.990 -2.985 25.290 4.170 ;
        RECT 25.625 -0.840 26.005 -0.460 ;
        RECT 26.330 -4.955 26.690 1.605 ;
        RECT 27.470 -0.205 27.795 1.660 ;
        RECT 28.135 -3.550 28.595 1.135 ;
        RECT 28.920 -1.005 29.370 7.815 ;
        RECT 31.105 0.820 31.535 3.810 ;
        RECT 28.850 -4.895 29.230 -4.515 ;
        RECT 31.740 -4.875 32.120 -3.500 ;
        RECT 32.510 -4.055 32.825 6.995 ;
        RECT 33.525 5.690 33.815 7.750 ;
        RECT 36.310 6.290 36.785 9.340 ;
        RECT 41.265 6.200 41.675 9.295 ;
        RECT 33.445 -2.165 33.770 0.205 ;
        RECT 35.095 -0.120 35.495 3.845 ;
        RECT 34.180 -5.905 34.525 -3.445 ;
        RECT 35.815 -4.225 36.140 -1.460 ;
        RECT 36.800 -2.190 37.205 1.140 ;
        RECT 41.450 -5.165 41.820 3.935 ;
        RECT 42.395 -4.100 42.685 7.735 ;
        RECT 45.845 6.175 46.255 9.270 ;
        RECT 50.300 5.630 50.610 8.145 ;
        RECT 46.210 -2.135 46.650 1.140 ;
        RECT 48.590 -0.120 49.115 3.820 ;
        RECT 47.750 -4.225 48.075 -1.460 ;
        RECT 50.265 -2.130 50.680 0.260 ;
        RECT 51.295 -3.570 51.610 7.115 ;
        RECT 52.625 0.820 53.110 3.830 ;
        RECT 51.995 -4.960 52.330 -3.610 ;
        RECT -7.795 -21.115 -7.380 -7.390 ;
        RECT 55.520 -8.170 56.075 2.845 ;
        RECT -6.355 -20.090 -5.940 -8.725 ;
        RECT 57.235 -9.590 57.705 -0.245 ;
        RECT 62.530 -9.400 63.055 2.020 ;
        RECT 64.660 -7.995 65.125 3.345 ;
        RECT 68.480 -4.045 68.835 7.040 ;
        RECT 72.225 5.680 72.515 7.740 ;
        RECT 74.995 6.280 75.495 9.330 ;
        RECT 79.965 6.190 80.375 9.285 ;
        RECT 79.005 4.530 79.315 4.560 ;
        RECT 69.805 0.810 70.275 3.800 ;
        RECT 72.155 -2.175 72.470 0.195 ;
        RECT 73.775 -0.130 74.195 3.835 ;
        RECT 70.440 -4.885 70.820 -3.510 ;
        RECT 72.880 -5.915 73.225 -3.455 ;
        RECT 74.515 -4.235 74.840 -1.470 ;
        RECT 75.500 -2.200 75.905 1.130 ;
        RECT 79.005 -1.570 79.320 4.530 ;
        RECT 80.150 -5.175 80.520 3.925 ;
        RECT 81.095 -4.110 81.385 7.725 ;
        RECT 84.545 6.165 84.955 9.260 ;
        RECT 89.000 5.620 89.310 8.135 ;
        RECT 93.250 7.320 93.630 7.700 ;
        RECT 95.380 7.320 95.760 7.700 ;
        RECT 81.990 -1.615 82.320 4.580 ;
        RECT 84.895 -2.145 85.350 1.130 ;
        RECT 87.255 -0.130 87.800 3.810 ;
        RECT 91.310 0.810 91.745 3.820 ;
        RECT 86.450 -4.235 86.775 -1.470 ;
        RECT 88.965 -2.140 89.380 0.250 ;
        RECT 92.505 -3.565 92.835 7.130 ;
        RECT 93.940 0.770 94.325 6.555 ;
        RECT 90.695 -4.970 91.030 -3.620 ;
        RECT 94.300 -3.985 94.725 0.290 ;
        RECT 96.000 -2.220 96.300 4.820 ;
        RECT 97.120 -2.825 97.420 4.105 ;
        RECT 98.430 -2.225 98.730 4.125 ;
        RECT 92.960 -4.895 93.340 -4.515 ;
        RECT 95.155 -4.910 95.535 -4.530 ;
        RECT 99.025 -4.970 99.315 4.810 ;
        RECT 99.745 -2.195 100.040 4.630 ;
        RECT 100.875 -2.735 101.175 4.075 ;
        RECT 101.665 -2.140 101.975 7.900 ;
        RECT 110.855 6.145 111.235 6.525 ;
        RECT 102.460 -2.210 102.760 4.620 ;
        RECT 103.585 -2.825 103.885 4.115 ;
        RECT 105.035 -2.950 105.315 0.085 ;
        RECT 105.795 -2.250 106.075 4.110 ;
        RECT 106.645 -2.250 106.945 4.570 ;
        RECT 107.785 -2.995 108.085 4.160 ;
        RECT 108.430 1.195 108.810 1.575 ;
        RECT 108.430 -0.860 108.810 -0.480 ;
        RECT 110.280 -0.980 110.595 3.345 ;
        RECT 110.890 1.095 111.170 2.625 ;
        RECT 111.460 -2.220 111.760 4.820 ;
        RECT 113.235 -1.465 113.535 2.595 ;
        RECT 110.755 -4.030 111.135 -3.650 ;
        RECT 114.485 -4.435 114.775 4.810 ;
        RECT 116.335 -2.735 116.635 4.075 ;
        RECT 117.125 -2.140 117.435 6.595 ;
        RECT 117.920 -2.210 118.220 4.620 ;
        RECT 119.725 -1.480 120.005 2.610 ;
        RECT 120.495 -2.950 120.775 0.085 ;
        RECT 123.245 -2.995 123.545 4.160 ;
        RECT 125.170 2.925 125.545 10.765 ;
        RECT 127.025 2.175 127.325 12.715 ;
        RECT -0.985 -22.610 -0.685 -15.680 ;
        RECT 0.325 -22.010 0.625 -15.660 ;
        RECT 1.640 -21.980 1.935 -15.155 ;
        RECT 5.480 -22.610 5.780 -15.670 ;
        RECT 7.690 -22.035 7.995 -15.675 ;
        RECT 8.540 -22.035 8.840 -15.215 ;
        RECT 10.350 -18.590 10.730 -18.210 ;
        RECT 12.135 -20.010 12.455 -17.880 ;
        RECT 10.565 -23.300 10.945 -20.280 ;
        RECT 12.745 -20.850 13.025 -18.445 ;
        RECT 13.355 -22.005 13.655 -14.965 ;
        RECT 14.475 -22.610 14.775 -15.680 ;
        RECT 15.785 -22.010 16.085 -15.660 ;
        RECT 16.380 -20.135 16.705 -14.975 ;
        RECT 17.100 -21.980 17.395 -15.155 ;
        RECT 18.230 -22.520 18.530 -15.710 ;
        RECT 19.020 -21.925 19.330 -15.735 ;
        RECT 19.815 -21.995 20.115 -15.165 ;
        RECT 20.940 -22.610 21.240 -15.670 ;
        RECT 22.390 -22.735 22.670 -19.700 ;
        RECT 23.150 -22.035 23.470 -15.675 ;
        RECT 24.000 -22.035 24.300 -15.215 ;
        RECT 25.140 -22.780 25.440 -15.625 ;
        RECT 25.775 -20.635 26.155 -20.255 ;
        RECT 26.480 -24.750 26.840 -18.190 ;
        RECT 27.620 -20.000 27.945 -18.135 ;
        RECT 28.285 -23.345 28.745 -18.660 ;
        RECT 29.070 -20.800 29.520 -11.980 ;
        RECT 31.255 -18.975 31.685 -15.985 ;
        RECT 29.000 -24.690 29.380 -24.310 ;
        RECT 31.890 -24.670 32.270 -23.295 ;
        RECT 32.660 -23.850 32.975 -12.800 ;
        RECT 33.675 -14.105 33.965 -12.045 ;
        RECT 36.460 -13.505 36.935 -10.455 ;
        RECT 41.415 -13.595 41.825 -10.500 ;
        RECT 33.595 -21.960 33.920 -19.590 ;
        RECT 35.245 -19.915 35.645 -15.950 ;
        RECT 34.330 -25.700 34.675 -23.240 ;
        RECT 35.965 -24.020 36.290 -21.255 ;
        RECT 36.950 -21.985 37.355 -18.655 ;
        RECT 41.600 -24.960 41.970 -15.860 ;
        RECT 42.545 -23.895 42.835 -12.060 ;
        RECT 45.995 -13.620 46.405 -10.525 ;
        RECT 50.450 -14.165 50.760 -11.650 ;
        RECT 46.360 -21.930 46.800 -18.655 ;
        RECT 48.740 -19.915 49.265 -15.975 ;
        RECT 47.900 -24.020 48.225 -21.255 ;
        RECT 50.415 -21.925 50.830 -19.535 ;
        RECT 51.445 -23.365 51.760 -12.680 ;
        RECT 52.775 -18.975 53.260 -15.965 ;
        RECT 52.145 -24.755 52.480 -23.405 ;
        RECT -8.140 -40.580 -7.785 -26.790 ;
        RECT 55.205 -27.420 55.655 -17.155 ;
        RECT -6.515 -39.725 -6.155 -28.390 ;
        RECT 56.370 -28.960 56.855 -20.075 ;
        RECT 62.675 -29.335 63.080 -17.805 ;
        RECT 64.750 -27.435 65.140 -16.335 ;
        RECT 68.520 -23.885 68.875 -12.800 ;
        RECT 72.265 -14.160 72.555 -12.100 ;
        RECT 75.035 -13.560 75.535 -10.510 ;
        RECT 80.005 -13.650 80.415 -10.555 ;
        RECT 79.045 -15.310 79.355 -15.280 ;
        RECT 69.845 -19.030 70.315 -16.040 ;
        RECT 72.195 -22.015 72.510 -19.645 ;
        RECT 73.815 -19.970 74.235 -16.005 ;
        RECT 70.480 -24.725 70.860 -23.350 ;
        RECT 72.920 -25.755 73.265 -23.295 ;
        RECT 74.555 -24.075 74.880 -21.310 ;
        RECT 75.540 -22.040 75.945 -18.710 ;
        RECT 79.045 -21.410 79.360 -15.310 ;
        RECT 80.190 -25.015 80.560 -15.915 ;
        RECT 81.135 -23.950 81.425 -12.115 ;
        RECT 84.585 -13.675 84.995 -10.580 ;
        RECT 89.040 -14.220 89.350 -11.705 ;
        RECT 93.290 -12.520 93.670 -12.140 ;
        RECT 95.420 -12.520 95.800 -12.140 ;
        RECT 82.030 -21.455 82.360 -15.260 ;
        RECT 84.935 -21.985 85.390 -18.710 ;
        RECT 87.295 -19.970 87.840 -16.030 ;
        RECT 91.350 -19.030 91.785 -16.020 ;
        RECT 86.490 -24.075 86.815 -21.310 ;
        RECT 89.005 -21.980 89.420 -19.590 ;
        RECT 92.545 -23.405 92.875 -12.710 ;
        RECT 93.980 -19.070 94.365 -13.285 ;
        RECT 90.735 -24.810 91.070 -23.460 ;
        RECT 94.340 -23.825 94.765 -19.550 ;
        RECT 96.040 -22.060 96.340 -15.020 ;
        RECT 97.160 -22.665 97.460 -15.735 ;
        RECT 98.470 -22.065 98.770 -15.715 ;
        RECT 93.000 -24.735 93.380 -24.355 ;
        RECT 95.195 -24.750 95.575 -24.370 ;
        RECT 99.065 -24.810 99.355 -15.030 ;
        RECT 99.785 -22.035 100.080 -15.210 ;
        RECT 100.915 -22.575 101.215 -15.765 ;
        RECT 101.705 -21.980 102.015 -11.940 ;
        RECT 110.895 -13.695 111.275 -13.315 ;
        RECT 102.500 -22.050 102.800 -15.220 ;
        RECT 103.625 -22.665 103.925 -15.725 ;
        RECT 105.075 -22.790 105.355 -19.755 ;
        RECT 105.835 -22.090 106.115 -15.730 ;
        RECT 106.685 -22.090 106.985 -15.270 ;
        RECT 107.825 -22.835 108.125 -15.680 ;
        RECT 108.470 -18.645 108.850 -18.265 ;
        RECT 108.470 -20.700 108.850 -20.320 ;
        RECT 110.320 -20.820 110.635 -16.495 ;
        RECT 110.930 -18.745 111.210 -17.215 ;
        RECT 111.500 -22.060 111.800 -15.020 ;
        RECT 113.275 -21.305 113.575 -17.245 ;
        RECT 110.795 -23.870 111.175 -23.490 ;
        RECT 114.525 -24.275 114.815 -15.030 ;
        RECT 116.375 -22.575 116.675 -15.765 ;
        RECT 117.165 -21.980 117.475 -13.245 ;
        RECT 117.960 -22.050 118.260 -15.220 ;
        RECT 119.765 -21.320 120.045 -17.230 ;
        RECT 120.535 -22.790 120.815 -19.755 ;
        RECT 123.285 -22.835 123.585 -15.680 ;
        RECT 125.485 -17.050 125.885 -8.310 ;
        RECT 127.065 -17.830 127.460 -6.950 ;
        RECT -1.030 -42.300 -0.730 -35.370 ;
        RECT 0.280 -41.700 0.580 -35.350 ;
        RECT 1.595 -41.670 1.890 -34.845 ;
        RECT 5.435 -42.300 5.735 -35.360 ;
        RECT 7.645 -41.725 7.950 -35.365 ;
        RECT 8.495 -41.725 8.795 -34.905 ;
        RECT 10.305 -38.280 10.685 -37.900 ;
        RECT 12.090 -39.700 12.410 -37.570 ;
        RECT 10.520 -42.990 10.900 -39.970 ;
        RECT 12.700 -40.540 12.980 -38.135 ;
        RECT 13.310 -41.695 13.610 -34.655 ;
        RECT 14.430 -42.300 14.730 -35.370 ;
        RECT 15.740 -41.700 16.040 -35.350 ;
        RECT 16.335 -39.825 16.660 -34.665 ;
        RECT 17.055 -41.670 17.350 -34.845 ;
        RECT 18.185 -42.210 18.485 -35.400 ;
        RECT 18.975 -41.615 19.285 -35.425 ;
        RECT 19.770 -41.685 20.070 -34.855 ;
        RECT 20.895 -42.300 21.195 -35.360 ;
        RECT 22.345 -42.425 22.625 -39.390 ;
        RECT 23.105 -41.725 23.425 -35.365 ;
        RECT 23.955 -41.725 24.255 -34.905 ;
        RECT 25.095 -42.470 25.395 -35.315 ;
        RECT 25.730 -40.325 26.110 -39.945 ;
        RECT 26.435 -44.440 26.795 -37.880 ;
        RECT 27.575 -39.690 27.900 -37.825 ;
        RECT 28.240 -43.035 28.700 -38.350 ;
        RECT 29.025 -40.490 29.475 -31.670 ;
        RECT 31.210 -38.665 31.640 -35.675 ;
        RECT 28.955 -44.380 29.335 -44.000 ;
        RECT 31.845 -44.360 32.225 -42.985 ;
        RECT 32.615 -43.540 32.930 -32.490 ;
        RECT 33.630 -33.795 33.920 -31.735 ;
        RECT 36.415 -33.195 36.890 -30.145 ;
        RECT 41.370 -33.285 41.780 -30.190 ;
        RECT 33.550 -41.650 33.875 -39.280 ;
        RECT 35.200 -39.605 35.600 -35.640 ;
        RECT 34.285 -45.390 34.630 -42.930 ;
        RECT 35.920 -43.710 36.245 -40.945 ;
        RECT 36.905 -41.675 37.310 -38.345 ;
        RECT 41.555 -44.650 41.925 -35.550 ;
        RECT 42.500 -43.585 42.790 -31.750 ;
        RECT 45.950 -33.310 46.360 -30.215 ;
        RECT 50.405 -33.855 50.715 -31.340 ;
        RECT 46.315 -41.620 46.755 -38.345 ;
        RECT 48.695 -39.605 49.220 -35.665 ;
        RECT 47.855 -43.710 48.180 -40.945 ;
        RECT 50.370 -41.615 50.785 -39.225 ;
        RECT 51.400 -43.055 51.715 -32.370 ;
        RECT 52.730 -38.665 53.215 -35.655 ;
        RECT 52.100 -44.445 52.435 -43.095 ;
        RECT -8.140 -60.345 -7.785 -46.290 ;
        RECT 55.205 -46.920 55.655 -36.805 ;
        RECT -6.515 -59.540 -6.155 -47.890 ;
        RECT 56.370 -48.460 56.855 -39.705 ;
        RECT 62.975 -49.085 63.380 -37.555 ;
        RECT 65.050 -47.185 65.440 -36.085 ;
        RECT 68.320 -43.610 68.675 -32.525 ;
        RECT 72.065 -33.885 72.355 -31.825 ;
        RECT 74.835 -33.285 75.335 -30.235 ;
        RECT 79.805 -33.375 80.215 -30.280 ;
        RECT 78.845 -35.035 79.155 -35.005 ;
        RECT 69.645 -38.755 70.115 -35.765 ;
        RECT 71.995 -41.740 72.310 -39.370 ;
        RECT 73.615 -39.695 74.035 -35.730 ;
        RECT 70.280 -44.450 70.660 -43.075 ;
        RECT 72.720 -45.480 73.065 -43.020 ;
        RECT 74.355 -43.800 74.680 -41.035 ;
        RECT 75.340 -41.765 75.745 -38.435 ;
        RECT 78.845 -41.135 79.160 -35.035 ;
        RECT 79.990 -44.740 80.360 -35.640 ;
        RECT 80.935 -43.675 81.225 -31.840 ;
        RECT 84.385 -33.400 84.795 -30.305 ;
        RECT 88.840 -33.945 89.150 -31.430 ;
        RECT 93.090 -32.245 93.470 -31.865 ;
        RECT 95.220 -32.245 95.600 -31.865 ;
        RECT 81.830 -41.180 82.160 -34.985 ;
        RECT 84.735 -41.710 85.190 -38.435 ;
        RECT 87.095 -39.695 87.640 -35.755 ;
        RECT 91.150 -38.755 91.585 -35.745 ;
        RECT 86.290 -43.800 86.615 -41.035 ;
        RECT 88.805 -41.705 89.220 -39.315 ;
        RECT 92.345 -43.130 92.675 -32.435 ;
        RECT 93.780 -38.795 94.165 -33.010 ;
        RECT 90.535 -44.535 90.870 -43.185 ;
        RECT 94.140 -43.550 94.565 -39.275 ;
        RECT 95.840 -41.785 96.140 -34.745 ;
        RECT 96.960 -42.390 97.260 -35.460 ;
        RECT 98.270 -41.790 98.570 -35.440 ;
        RECT 92.800 -44.460 93.180 -44.080 ;
        RECT 94.995 -44.475 95.375 -44.095 ;
        RECT 98.865 -44.535 99.155 -34.755 ;
        RECT 99.585 -41.760 99.880 -34.935 ;
        RECT 100.715 -42.300 101.015 -35.490 ;
        RECT 101.505 -41.705 101.815 -31.665 ;
        RECT 110.695 -33.420 111.075 -33.040 ;
        RECT 102.300 -41.775 102.600 -34.945 ;
        RECT 103.425 -42.390 103.725 -35.450 ;
        RECT 104.875 -42.515 105.155 -39.480 ;
        RECT 105.635 -41.815 105.915 -35.455 ;
        RECT 106.485 -41.815 106.785 -34.995 ;
        RECT 107.625 -42.560 107.925 -35.405 ;
        RECT 108.270 -38.370 108.650 -37.990 ;
        RECT 108.270 -40.425 108.650 -40.045 ;
        RECT 110.120 -40.545 110.435 -36.220 ;
        RECT 110.730 -38.470 111.010 -36.940 ;
        RECT 111.300 -41.785 111.600 -34.745 ;
        RECT 113.075 -41.030 113.375 -36.970 ;
        RECT 110.595 -43.595 110.975 -43.215 ;
        RECT 114.325 -44.000 114.615 -34.755 ;
        RECT 116.175 -42.300 116.475 -35.490 ;
        RECT 116.965 -41.705 117.275 -32.970 ;
        RECT 117.760 -41.775 118.060 -34.945 ;
        RECT 119.565 -41.045 119.845 -36.955 ;
        RECT 120.335 -42.515 120.615 -39.480 ;
        RECT 123.085 -42.560 123.385 -35.405 ;
        RECT 125.125 -36.665 125.500 -28.465 ;
        RECT 126.870 -37.470 127.170 -26.475 ;
        RECT -0.840 -62.010 -0.540 -55.080 ;
        RECT 0.470 -61.410 0.770 -55.060 ;
        RECT 1.785 -61.380 2.080 -54.555 ;
        RECT 5.625 -62.010 5.925 -55.070 ;
        RECT 7.835 -61.435 8.140 -55.075 ;
        RECT 8.685 -61.435 8.985 -54.615 ;
        RECT 10.495 -57.990 10.875 -57.610 ;
        RECT 12.280 -59.410 12.600 -57.280 ;
        RECT 10.710 -62.700 11.090 -59.680 ;
        RECT 12.890 -60.250 13.170 -57.845 ;
        RECT 13.500 -61.405 13.800 -54.365 ;
        RECT 14.620 -62.010 14.920 -55.080 ;
        RECT 15.930 -61.410 16.230 -55.060 ;
        RECT 16.525 -59.535 16.850 -54.375 ;
        RECT 17.245 -61.380 17.540 -54.555 ;
        RECT 18.375 -61.920 18.675 -55.110 ;
        RECT 19.165 -61.325 19.475 -55.135 ;
        RECT 19.960 -61.395 20.260 -54.565 ;
        RECT 21.085 -62.010 21.385 -55.070 ;
        RECT 22.535 -62.135 22.815 -59.100 ;
        RECT 23.295 -61.435 23.615 -55.075 ;
        RECT 24.145 -61.435 24.445 -54.615 ;
        RECT 25.285 -62.180 25.585 -55.025 ;
        RECT 25.920 -60.035 26.300 -59.655 ;
        RECT 26.625 -64.150 26.985 -57.590 ;
        RECT 27.765 -59.400 28.090 -57.535 ;
        RECT 28.430 -62.745 28.890 -58.060 ;
        RECT 29.215 -60.200 29.665 -51.380 ;
        RECT 31.400 -58.375 31.830 -55.385 ;
        RECT 29.145 -64.090 29.525 -63.710 ;
        RECT 32.035 -64.070 32.415 -62.695 ;
        RECT 32.805 -63.250 33.120 -52.200 ;
        RECT 33.820 -53.505 34.110 -51.445 ;
        RECT 36.605 -52.905 37.080 -49.855 ;
        RECT 41.560 -52.995 41.970 -49.900 ;
        RECT 33.740 -61.360 34.065 -58.990 ;
        RECT 35.390 -59.315 35.790 -55.350 ;
        RECT 34.475 -65.100 34.820 -62.640 ;
        RECT 36.110 -63.420 36.435 -60.655 ;
        RECT 37.095 -61.385 37.500 -58.055 ;
        RECT 41.745 -64.360 42.115 -55.260 ;
        RECT 42.690 -63.295 42.980 -51.460 ;
        RECT 46.140 -53.020 46.550 -49.925 ;
        RECT 50.595 -53.565 50.905 -51.050 ;
        RECT 46.505 -61.330 46.945 -58.055 ;
        RECT 48.885 -59.315 49.410 -55.375 ;
        RECT 48.045 -63.420 48.370 -60.655 ;
        RECT 50.560 -61.325 50.975 -58.935 ;
        RECT 51.590 -62.765 51.905 -52.080 ;
        RECT 52.920 -58.375 53.405 -55.365 ;
        RECT 52.290 -64.155 52.625 -62.805 ;
        RECT -7.930 -80.120 -7.575 -66.330 ;
        RECT 55.415 -66.960 55.865 -56.460 ;
        RECT -6.305 -79.265 -5.945 -67.930 ;
        RECT 56.580 -68.500 57.065 -59.260 ;
        RECT 62.995 -68.745 63.400 -57.215 ;
        RECT 65.070 -66.845 65.460 -55.745 ;
        RECT 68.475 -63.255 68.830 -52.170 ;
        RECT 72.220 -53.530 72.510 -51.470 ;
        RECT 74.990 -52.930 75.490 -49.880 ;
        RECT 79.960 -53.020 80.370 -49.925 ;
        RECT 79.000 -54.680 79.310 -54.650 ;
        RECT 69.800 -58.400 70.270 -55.410 ;
        RECT 72.150 -61.385 72.465 -59.015 ;
        RECT 73.770 -59.340 74.190 -55.375 ;
        RECT 70.435 -64.095 70.815 -62.720 ;
        RECT 72.875 -65.125 73.220 -62.665 ;
        RECT 74.510 -63.445 74.835 -60.680 ;
        RECT 75.495 -61.410 75.900 -58.080 ;
        RECT 79.000 -60.780 79.315 -54.680 ;
        RECT 80.145 -64.385 80.515 -55.285 ;
        RECT 81.090 -63.320 81.380 -51.485 ;
        RECT 84.540 -53.045 84.950 -49.950 ;
        RECT 88.995 -53.590 89.305 -51.075 ;
        RECT 93.245 -51.890 93.625 -51.510 ;
        RECT 95.375 -51.890 95.755 -51.510 ;
        RECT 81.985 -60.825 82.315 -54.630 ;
        RECT 84.890 -61.355 85.345 -58.080 ;
        RECT 87.250 -59.340 87.795 -55.400 ;
        RECT 91.305 -58.400 91.740 -55.390 ;
        RECT 86.445 -63.445 86.770 -60.680 ;
        RECT 88.960 -61.350 89.375 -58.960 ;
        RECT 92.500 -62.775 92.830 -52.080 ;
        RECT 93.935 -58.440 94.320 -52.655 ;
        RECT 90.690 -64.180 91.025 -62.830 ;
        RECT 94.295 -63.195 94.720 -58.920 ;
        RECT 95.995 -61.430 96.295 -54.390 ;
        RECT 97.115 -62.035 97.415 -55.105 ;
        RECT 98.425 -61.435 98.725 -55.085 ;
        RECT 92.955 -64.105 93.335 -63.725 ;
        RECT 95.150 -64.120 95.530 -63.740 ;
        RECT 99.020 -64.180 99.310 -54.400 ;
        RECT 99.740 -61.405 100.035 -54.580 ;
        RECT 100.870 -61.945 101.170 -55.135 ;
        RECT 101.660 -61.350 101.970 -51.310 ;
        RECT 110.850 -53.065 111.230 -52.685 ;
        RECT 102.455 -61.420 102.755 -54.590 ;
        RECT 103.580 -62.035 103.880 -55.095 ;
        RECT 105.030 -62.160 105.310 -59.125 ;
        RECT 105.790 -61.460 106.070 -55.100 ;
        RECT 106.640 -61.460 106.940 -54.640 ;
        RECT 107.780 -62.205 108.080 -55.050 ;
        RECT 108.425 -58.015 108.805 -57.635 ;
        RECT 108.425 -60.070 108.805 -59.690 ;
        RECT 110.275 -60.190 110.590 -55.865 ;
        RECT 110.885 -58.115 111.165 -56.585 ;
        RECT 111.455 -61.430 111.755 -54.390 ;
        RECT 113.230 -60.675 113.530 -56.615 ;
        RECT 110.750 -63.240 111.130 -62.860 ;
        RECT 114.480 -63.645 114.770 -54.400 ;
        RECT 116.330 -61.945 116.630 -55.135 ;
        RECT 117.120 -61.350 117.430 -52.615 ;
        RECT 117.915 -61.420 118.215 -54.590 ;
        RECT 119.720 -60.690 120.000 -56.600 ;
        RECT 120.490 -62.160 120.770 -59.125 ;
        RECT 123.240 -62.205 123.540 -55.050 ;
        RECT 125.425 -56.415 125.800 -48.215 ;
        RECT 127.170 -57.220 127.470 -46.225 ;
        RECT -1.035 -81.850 -0.735 -74.920 ;
        RECT 0.275 -81.250 0.575 -74.900 ;
        RECT 1.590 -81.220 1.885 -74.395 ;
        RECT 5.430 -81.850 5.730 -74.910 ;
        RECT 7.640 -81.275 7.945 -74.915 ;
        RECT 8.490 -81.275 8.790 -74.455 ;
        RECT 10.300 -77.830 10.680 -77.450 ;
        RECT 12.085 -79.250 12.405 -77.120 ;
        RECT 10.515 -82.540 10.895 -79.520 ;
        RECT 12.695 -80.090 12.975 -77.685 ;
        RECT 13.305 -81.245 13.605 -74.205 ;
        RECT 14.425 -81.850 14.725 -74.920 ;
        RECT 15.735 -81.250 16.035 -74.900 ;
        RECT 16.330 -79.375 16.655 -74.215 ;
        RECT 17.050 -81.220 17.345 -74.395 ;
        RECT 18.180 -81.760 18.480 -74.950 ;
        RECT 18.970 -81.165 19.280 -74.975 ;
        RECT 19.765 -81.235 20.065 -74.405 ;
        RECT 20.890 -81.850 21.190 -74.910 ;
        RECT 22.340 -81.975 22.620 -78.940 ;
        RECT 23.100 -81.275 23.420 -74.915 ;
        RECT 23.950 -81.275 24.250 -74.455 ;
        RECT 25.090 -82.020 25.390 -74.865 ;
        RECT 25.725 -79.875 26.105 -79.495 ;
        RECT 26.430 -83.990 26.790 -77.430 ;
        RECT 27.570 -79.240 27.895 -77.375 ;
        RECT 28.235 -82.585 28.695 -77.900 ;
        RECT 29.020 -80.040 29.470 -71.220 ;
        RECT 31.205 -78.215 31.635 -75.225 ;
        RECT 28.950 -83.930 29.330 -83.550 ;
        RECT 31.840 -83.910 32.220 -82.535 ;
        RECT 32.610 -83.090 32.925 -72.040 ;
        RECT 33.625 -73.345 33.915 -71.285 ;
        RECT 36.410 -72.745 36.885 -69.695 ;
        RECT 41.365 -72.835 41.775 -69.740 ;
        RECT 33.545 -81.200 33.870 -78.830 ;
        RECT 35.195 -79.155 35.595 -75.190 ;
        RECT 34.280 -84.940 34.625 -82.480 ;
        RECT 35.915 -83.260 36.240 -80.495 ;
        RECT 36.900 -81.225 37.305 -77.895 ;
        RECT 41.550 -84.200 41.920 -75.100 ;
        RECT 42.495 -83.135 42.785 -71.300 ;
        RECT 45.945 -72.860 46.355 -69.765 ;
        RECT 50.400 -73.405 50.710 -70.890 ;
        RECT 46.310 -81.170 46.750 -77.895 ;
        RECT 48.690 -79.155 49.215 -75.215 ;
        RECT 47.850 -83.260 48.175 -80.495 ;
        RECT 50.365 -81.165 50.780 -78.775 ;
        RECT 51.395 -82.605 51.710 -71.920 ;
        RECT 52.725 -78.215 53.210 -75.205 ;
        RECT 52.095 -83.995 52.430 -82.645 ;
        RECT -7.975 -99.910 -7.620 -86.120 ;
        RECT 55.370 -86.750 55.820 -76.260 ;
        RECT -6.350 -99.005 -5.990 -87.720 ;
        RECT 56.535 -88.290 57.020 -79.130 ;
        RECT 62.995 -88.480 63.400 -76.950 ;
        RECT 65.070 -86.580 65.460 -75.480 ;
        RECT 68.475 -83.050 68.830 -71.965 ;
        RECT 72.220 -73.325 72.510 -71.265 ;
        RECT 74.990 -72.725 75.490 -69.675 ;
        RECT 79.960 -72.815 80.370 -69.720 ;
        RECT 79.000 -74.475 79.310 -74.445 ;
        RECT 69.800 -78.195 70.270 -75.205 ;
        RECT 72.150 -81.180 72.465 -78.810 ;
        RECT 73.770 -79.135 74.190 -75.170 ;
        RECT 70.435 -83.890 70.815 -82.515 ;
        RECT 72.875 -84.920 73.220 -82.460 ;
        RECT 74.510 -83.240 74.835 -80.475 ;
        RECT 75.495 -81.205 75.900 -77.875 ;
        RECT 79.000 -80.575 79.315 -74.475 ;
        RECT 80.145 -84.180 80.515 -75.080 ;
        RECT 81.090 -83.115 81.380 -71.280 ;
        RECT 84.540 -72.840 84.950 -69.745 ;
        RECT 88.995 -73.385 89.305 -70.870 ;
        RECT 93.245 -71.685 93.625 -71.305 ;
        RECT 95.375 -71.685 95.755 -71.305 ;
        RECT 81.985 -80.620 82.315 -74.425 ;
        RECT 84.890 -81.150 85.345 -77.875 ;
        RECT 87.250 -79.135 87.795 -75.195 ;
        RECT 91.305 -78.195 91.740 -75.185 ;
        RECT 86.445 -83.240 86.770 -80.475 ;
        RECT 88.960 -81.145 89.375 -78.755 ;
        RECT 92.500 -82.570 92.830 -71.875 ;
        RECT 93.935 -78.235 94.320 -72.450 ;
        RECT 90.690 -83.975 91.025 -82.625 ;
        RECT 94.295 -82.990 94.720 -78.715 ;
        RECT 95.995 -81.225 96.295 -74.185 ;
        RECT 97.115 -81.830 97.415 -74.900 ;
        RECT 98.425 -81.230 98.725 -74.880 ;
        RECT 92.955 -83.900 93.335 -83.520 ;
        RECT 95.150 -83.915 95.530 -83.535 ;
        RECT 99.020 -83.975 99.310 -74.195 ;
        RECT 99.740 -81.200 100.035 -74.375 ;
        RECT 100.870 -81.740 101.170 -74.930 ;
        RECT 101.660 -81.145 101.970 -71.105 ;
        RECT 110.850 -72.860 111.230 -72.480 ;
        RECT 102.455 -81.215 102.755 -74.385 ;
        RECT 103.580 -81.830 103.880 -74.890 ;
        RECT 105.030 -81.955 105.310 -78.920 ;
        RECT 105.790 -81.255 106.070 -74.895 ;
        RECT 106.640 -81.255 106.940 -74.435 ;
        RECT 107.780 -82.000 108.080 -74.845 ;
        RECT 108.425 -77.810 108.805 -77.430 ;
        RECT 108.425 -79.865 108.805 -79.485 ;
        RECT 110.275 -79.985 110.590 -75.660 ;
        RECT 110.885 -77.910 111.165 -76.380 ;
        RECT 111.455 -81.225 111.755 -74.185 ;
        RECT 113.230 -80.470 113.530 -76.410 ;
        RECT 110.750 -83.035 111.130 -82.655 ;
        RECT 114.480 -83.440 114.770 -74.195 ;
        RECT 116.330 -81.740 116.630 -74.930 ;
        RECT 117.120 -81.145 117.430 -72.410 ;
        RECT 117.915 -81.215 118.215 -74.385 ;
        RECT 119.720 -80.485 120.000 -76.395 ;
        RECT 120.490 -81.955 120.770 -78.920 ;
        RECT 123.240 -82.000 123.540 -74.845 ;
        RECT 125.445 -76.075 125.820 -67.875 ;
        RECT 127.190 -76.880 127.490 -65.885 ;
        RECT -1.165 -101.560 -0.865 -94.630 ;
        RECT 0.145 -100.960 0.445 -94.610 ;
        RECT 1.460 -100.930 1.755 -94.105 ;
        RECT 5.300 -101.560 5.600 -94.620 ;
        RECT 7.510 -100.985 7.815 -94.625 ;
        RECT 8.360 -100.985 8.660 -94.165 ;
        RECT 10.170 -97.540 10.550 -97.160 ;
        RECT 11.955 -98.960 12.275 -96.830 ;
        RECT 10.385 -102.250 10.765 -99.230 ;
        RECT 12.565 -99.800 12.845 -97.395 ;
        RECT 13.175 -100.955 13.475 -93.915 ;
        RECT 14.295 -101.560 14.595 -94.630 ;
        RECT 15.605 -100.960 15.905 -94.610 ;
        RECT 16.200 -99.085 16.525 -93.925 ;
        RECT 16.920 -100.930 17.215 -94.105 ;
        RECT 18.050 -101.470 18.350 -94.660 ;
        RECT 18.840 -100.875 19.150 -94.685 ;
        RECT 19.635 -100.945 19.935 -94.115 ;
        RECT 20.760 -101.560 21.060 -94.620 ;
        RECT 22.210 -101.685 22.490 -98.650 ;
        RECT 22.970 -100.985 23.290 -94.625 ;
        RECT 23.820 -100.985 24.120 -94.165 ;
        RECT 24.960 -101.730 25.260 -94.575 ;
        RECT 25.595 -99.585 25.975 -99.205 ;
        RECT 26.300 -103.700 26.660 -97.140 ;
        RECT 27.440 -98.950 27.765 -97.085 ;
        RECT 28.105 -102.295 28.565 -97.610 ;
        RECT 28.890 -99.750 29.340 -90.930 ;
        RECT 31.075 -97.925 31.505 -94.935 ;
        RECT 28.820 -103.640 29.200 -103.260 ;
        RECT 31.710 -103.620 32.090 -102.245 ;
        RECT 32.480 -102.800 32.795 -91.750 ;
        RECT 33.495 -93.055 33.785 -90.995 ;
        RECT 36.280 -92.455 36.755 -89.405 ;
        RECT 41.235 -92.545 41.645 -89.450 ;
        RECT 33.415 -100.910 33.740 -98.540 ;
        RECT 35.065 -98.865 35.465 -94.900 ;
        RECT 34.150 -104.650 34.495 -102.190 ;
        RECT 35.785 -102.970 36.110 -100.205 ;
        RECT 36.770 -100.935 37.175 -97.605 ;
        RECT 41.420 -103.910 41.790 -94.810 ;
        RECT 42.365 -102.845 42.655 -91.010 ;
        RECT 45.815 -92.570 46.225 -89.475 ;
        RECT 50.270 -93.115 50.580 -90.600 ;
        RECT 46.180 -100.880 46.620 -97.605 ;
        RECT 48.560 -98.865 49.085 -94.925 ;
        RECT 47.720 -102.970 48.045 -100.205 ;
        RECT 50.235 -100.875 50.650 -98.485 ;
        RECT 51.265 -102.315 51.580 -91.630 ;
        RECT 52.595 -97.925 53.080 -94.915 ;
        RECT 51.965 -103.705 52.300 -102.355 ;
        RECT -8.280 -119.670 -7.925 -105.750 ;
        RECT 55.065 -106.380 55.515 -96.115 ;
        RECT -6.655 -118.765 -6.295 -107.350 ;
        RECT 56.230 -107.920 56.715 -99.035 ;
        RECT 62.895 -108.185 63.300 -96.655 ;
        RECT 64.970 -106.285 65.360 -95.185 ;
        RECT 68.395 -102.805 68.750 -91.720 ;
        RECT 72.140 -93.080 72.430 -91.020 ;
        RECT 74.910 -92.480 75.410 -89.430 ;
        RECT 79.880 -92.570 80.290 -89.475 ;
        RECT 78.920 -94.230 79.230 -94.200 ;
        RECT 69.720 -97.950 70.190 -94.960 ;
        RECT 72.070 -100.935 72.385 -98.565 ;
        RECT 73.690 -98.890 74.110 -94.925 ;
        RECT 70.355 -103.645 70.735 -102.270 ;
        RECT 72.795 -104.675 73.140 -102.215 ;
        RECT 74.430 -102.995 74.755 -100.230 ;
        RECT 75.415 -100.960 75.820 -97.630 ;
        RECT 78.920 -100.330 79.235 -94.230 ;
        RECT 80.065 -103.935 80.435 -94.835 ;
        RECT 81.010 -102.870 81.300 -91.035 ;
        RECT 84.460 -92.595 84.870 -89.500 ;
        RECT 88.915 -93.140 89.225 -90.625 ;
        RECT 93.165 -91.440 93.545 -91.060 ;
        RECT 95.295 -91.440 95.675 -91.060 ;
        RECT 81.905 -100.375 82.235 -94.180 ;
        RECT 84.810 -100.905 85.265 -97.630 ;
        RECT 87.170 -98.890 87.715 -94.950 ;
        RECT 91.225 -97.950 91.660 -94.940 ;
        RECT 86.365 -102.995 86.690 -100.230 ;
        RECT 88.880 -100.900 89.295 -98.510 ;
        RECT 92.420 -102.325 92.750 -91.630 ;
        RECT 93.855 -97.990 94.240 -92.205 ;
        RECT 90.610 -103.730 90.945 -102.380 ;
        RECT 94.215 -102.745 94.640 -98.470 ;
        RECT 95.915 -100.980 96.215 -93.940 ;
        RECT 97.035 -101.585 97.335 -94.655 ;
        RECT 98.345 -100.985 98.645 -94.635 ;
        RECT 92.875 -103.655 93.255 -103.275 ;
        RECT 95.070 -103.670 95.450 -103.290 ;
        RECT 98.940 -103.730 99.230 -93.950 ;
        RECT 99.660 -100.955 99.955 -94.130 ;
        RECT 100.790 -101.495 101.090 -94.685 ;
        RECT 101.580 -100.900 101.890 -90.860 ;
        RECT 110.770 -92.615 111.150 -92.235 ;
        RECT 102.375 -100.970 102.675 -94.140 ;
        RECT 103.500 -101.585 103.800 -94.645 ;
        RECT 104.950 -101.710 105.230 -98.675 ;
        RECT 105.710 -101.010 105.990 -94.650 ;
        RECT 106.560 -101.010 106.860 -94.190 ;
        RECT 107.700 -101.755 108.000 -94.600 ;
        RECT 108.345 -97.565 108.725 -97.185 ;
        RECT 108.345 -99.620 108.725 -99.240 ;
        RECT 110.195 -99.740 110.510 -95.415 ;
        RECT 110.805 -97.665 111.085 -96.135 ;
        RECT 111.375 -100.980 111.675 -93.940 ;
        RECT 113.150 -100.225 113.450 -96.165 ;
        RECT 110.670 -102.790 111.050 -102.410 ;
        RECT 114.400 -103.195 114.690 -93.950 ;
        RECT 116.250 -101.495 116.550 -94.685 ;
        RECT 117.040 -100.900 117.350 -92.165 ;
        RECT 117.835 -100.970 118.135 -94.140 ;
        RECT 119.640 -100.240 119.920 -96.150 ;
        RECT 120.410 -101.710 120.690 -98.675 ;
        RECT 123.160 -101.755 123.460 -94.600 ;
        RECT 125.445 -95.895 125.820 -87.610 ;
        RECT 127.190 -96.615 127.490 -85.620 ;
        RECT -1.035 -121.320 -0.735 -114.390 ;
        RECT 0.275 -120.720 0.575 -114.370 ;
        RECT 1.590 -120.690 1.885 -113.865 ;
        RECT 5.430 -121.320 5.730 -114.380 ;
        RECT 7.640 -120.745 7.945 -114.385 ;
        RECT 8.490 -120.745 8.790 -113.925 ;
        RECT 10.300 -117.300 10.680 -116.920 ;
        RECT 12.085 -118.720 12.405 -116.590 ;
        RECT 10.515 -122.010 10.895 -118.990 ;
        RECT 12.695 -119.560 12.975 -117.155 ;
        RECT 13.305 -120.715 13.605 -113.675 ;
        RECT 14.425 -121.320 14.725 -114.390 ;
        RECT 15.735 -120.720 16.035 -114.370 ;
        RECT 16.330 -118.845 16.655 -113.685 ;
        RECT 17.050 -120.690 17.345 -113.865 ;
        RECT 18.180 -121.230 18.480 -114.420 ;
        RECT 18.970 -120.635 19.280 -114.445 ;
        RECT 19.765 -120.705 20.065 -113.875 ;
        RECT 20.890 -121.320 21.190 -114.380 ;
        RECT 22.340 -121.445 22.620 -118.410 ;
        RECT 23.100 -120.745 23.420 -114.385 ;
        RECT 23.950 -120.745 24.250 -113.925 ;
        RECT 25.090 -121.490 25.390 -114.335 ;
        RECT 25.725 -119.345 26.105 -118.965 ;
        RECT 26.430 -123.460 26.790 -116.900 ;
        RECT 27.570 -118.710 27.895 -116.845 ;
        RECT 28.235 -122.055 28.695 -117.370 ;
        RECT 29.020 -119.510 29.470 -110.690 ;
        RECT 31.205 -117.685 31.635 -114.695 ;
        RECT 28.950 -123.400 29.330 -123.020 ;
        RECT 31.840 -123.380 32.220 -122.005 ;
        RECT 32.610 -122.560 32.925 -111.510 ;
        RECT 33.625 -112.815 33.915 -110.755 ;
        RECT 36.410 -112.215 36.885 -109.165 ;
        RECT 41.365 -112.305 41.775 -109.210 ;
        RECT 33.545 -120.670 33.870 -118.300 ;
        RECT 35.195 -118.625 35.595 -114.660 ;
        RECT 34.280 -124.410 34.625 -121.950 ;
        RECT 35.915 -122.730 36.240 -119.965 ;
        RECT 36.900 -120.695 37.305 -117.365 ;
        RECT 41.550 -123.670 41.920 -114.570 ;
        RECT 42.495 -122.605 42.785 -110.770 ;
        RECT 45.945 -112.330 46.355 -109.235 ;
        RECT 50.400 -112.875 50.710 -110.360 ;
        RECT 46.310 -120.640 46.750 -117.365 ;
        RECT 48.690 -118.625 49.215 -114.685 ;
        RECT 47.850 -122.730 48.175 -119.965 ;
        RECT 50.365 -120.635 50.780 -118.245 ;
        RECT 51.395 -122.075 51.710 -111.390 ;
        RECT 52.725 -117.685 53.210 -114.675 ;
        RECT 52.095 -123.465 52.430 -122.115 ;
        RECT -8.185 -139.435 -7.830 -125.525 ;
        RECT 55.160 -126.155 55.610 -115.890 ;
        RECT -6.560 -138.515 -6.200 -127.125 ;
        RECT 56.325 -127.695 56.810 -118.810 ;
        RECT 63.155 -128.340 63.560 -116.460 ;
        RECT 65.230 -126.440 65.620 -114.860 ;
        RECT 68.500 -122.520 68.855 -111.435 ;
        RECT 72.245 -112.795 72.535 -110.735 ;
        RECT 75.015 -112.195 75.515 -109.145 ;
        RECT 79.985 -112.285 80.395 -109.190 ;
        RECT 79.025 -113.945 79.335 -113.915 ;
        RECT 69.825 -117.665 70.295 -114.675 ;
        RECT 72.175 -120.650 72.490 -118.280 ;
        RECT 73.795 -118.605 74.215 -114.640 ;
        RECT 70.460 -123.360 70.840 -121.985 ;
        RECT 72.900 -124.390 73.245 -121.930 ;
        RECT 74.535 -122.710 74.860 -119.945 ;
        RECT 75.520 -120.675 75.925 -117.345 ;
        RECT 79.025 -120.045 79.340 -113.945 ;
        RECT 80.170 -123.650 80.540 -114.550 ;
        RECT 81.115 -122.585 81.405 -110.750 ;
        RECT 84.565 -112.310 84.975 -109.215 ;
        RECT 89.020 -112.855 89.330 -110.340 ;
        RECT 93.270 -111.155 93.650 -110.775 ;
        RECT 95.400 -111.155 95.780 -110.775 ;
        RECT 82.010 -120.090 82.340 -113.895 ;
        RECT 84.915 -120.620 85.370 -117.345 ;
        RECT 87.275 -118.605 87.820 -114.665 ;
        RECT 91.330 -117.665 91.765 -114.655 ;
        RECT 86.470 -122.710 86.795 -119.945 ;
        RECT 88.985 -120.615 89.400 -118.225 ;
        RECT 92.525 -122.040 92.855 -111.345 ;
        RECT 93.960 -117.705 94.345 -111.920 ;
        RECT 90.715 -123.445 91.050 -122.095 ;
        RECT 94.320 -122.460 94.745 -118.185 ;
        RECT 96.020 -120.695 96.320 -113.655 ;
        RECT 97.140 -121.300 97.440 -114.370 ;
        RECT 98.450 -120.700 98.750 -114.350 ;
        RECT 92.980 -123.370 93.360 -122.990 ;
        RECT 95.175 -123.385 95.555 -123.005 ;
        RECT 99.045 -123.445 99.335 -113.665 ;
        RECT 99.765 -120.670 100.060 -113.845 ;
        RECT 100.895 -121.210 101.195 -114.400 ;
        RECT 101.685 -120.615 101.995 -110.575 ;
        RECT 110.875 -112.330 111.255 -111.950 ;
        RECT 102.480 -120.685 102.780 -113.855 ;
        RECT 103.605 -121.300 103.905 -114.360 ;
        RECT 105.055 -121.425 105.335 -118.390 ;
        RECT 105.815 -120.725 106.095 -114.365 ;
        RECT 106.665 -120.725 106.965 -113.905 ;
        RECT 107.805 -121.470 108.105 -114.315 ;
        RECT 108.450 -117.280 108.830 -116.900 ;
        RECT 108.450 -119.335 108.830 -118.955 ;
        RECT 110.300 -119.455 110.615 -115.130 ;
        RECT 110.910 -117.380 111.190 -115.850 ;
        RECT 111.480 -120.695 111.780 -113.655 ;
        RECT 113.255 -119.940 113.555 -115.880 ;
        RECT 110.775 -122.505 111.155 -122.125 ;
        RECT 114.505 -122.910 114.795 -113.665 ;
        RECT 116.355 -121.210 116.655 -114.400 ;
        RECT 117.145 -120.615 117.455 -111.880 ;
        RECT 117.940 -120.685 118.240 -113.855 ;
        RECT 119.745 -119.955 120.025 -115.865 ;
        RECT 120.515 -121.425 120.795 -118.390 ;
        RECT 123.265 -121.470 123.565 -114.315 ;
        RECT 125.345 -115.595 125.720 -107.315 ;
        RECT 127.090 -116.435 127.390 -105.325 ;
        RECT -1.085 -141.130 -0.785 -134.200 ;
        RECT 0.225 -140.530 0.525 -134.180 ;
        RECT 1.540 -140.500 1.835 -133.675 ;
        RECT 5.380 -141.130 5.680 -134.190 ;
        RECT 7.590 -140.555 7.895 -134.195 ;
        RECT 8.440 -140.555 8.740 -133.735 ;
        RECT 10.250 -137.110 10.630 -136.730 ;
        RECT 12.035 -138.530 12.355 -136.400 ;
        RECT 10.465 -141.820 10.845 -138.800 ;
        RECT 12.645 -139.370 12.925 -136.965 ;
        RECT 13.255 -140.525 13.555 -133.485 ;
        RECT 14.375 -141.130 14.675 -134.200 ;
        RECT 15.685 -140.530 15.985 -134.180 ;
        RECT 16.280 -138.655 16.605 -133.495 ;
        RECT 17.000 -140.500 17.295 -133.675 ;
        RECT 18.130 -141.040 18.430 -134.230 ;
        RECT 18.920 -140.445 19.230 -134.255 ;
        RECT 19.715 -140.515 20.015 -133.685 ;
        RECT 20.840 -141.130 21.140 -134.190 ;
        RECT 22.290 -141.255 22.570 -138.220 ;
        RECT 23.050 -140.555 23.370 -134.195 ;
        RECT 23.900 -140.555 24.200 -133.735 ;
        RECT 25.040 -141.300 25.340 -134.145 ;
        RECT 25.675 -139.155 26.055 -138.775 ;
        RECT 26.380 -143.270 26.740 -136.710 ;
        RECT 27.520 -138.520 27.845 -136.655 ;
        RECT 28.185 -141.865 28.645 -137.180 ;
        RECT 28.970 -139.320 29.420 -130.500 ;
        RECT 31.155 -137.495 31.585 -134.505 ;
        RECT 28.900 -143.210 29.280 -142.830 ;
        RECT 31.790 -143.190 32.170 -141.815 ;
        RECT 32.560 -142.370 32.875 -131.320 ;
        RECT 33.575 -132.625 33.865 -130.565 ;
        RECT 36.360 -132.025 36.835 -128.975 ;
        RECT 41.315 -132.115 41.725 -129.020 ;
        RECT 33.495 -140.480 33.820 -138.110 ;
        RECT 35.145 -138.435 35.545 -134.470 ;
        RECT 34.230 -144.220 34.575 -141.760 ;
        RECT 35.865 -142.540 36.190 -139.775 ;
        RECT 36.850 -140.505 37.255 -137.175 ;
        RECT 41.500 -143.480 41.870 -134.380 ;
        RECT 42.445 -142.415 42.735 -130.580 ;
        RECT 45.895 -132.140 46.305 -129.045 ;
        RECT 50.350 -132.685 50.660 -130.170 ;
        RECT 46.260 -140.450 46.700 -137.175 ;
        RECT 48.640 -138.435 49.165 -134.495 ;
        RECT 47.800 -142.540 48.125 -139.775 ;
        RECT 50.315 -140.445 50.730 -138.055 ;
        RECT 51.345 -141.885 51.660 -131.200 ;
        RECT 52.675 -137.495 53.160 -134.485 ;
        RECT 52.045 -143.275 52.380 -141.925 ;
        RECT -8.185 -159.275 -7.830 -145.335 ;
        RECT 55.160 -145.965 55.610 -135.700 ;
        RECT -6.560 -158.485 -6.200 -146.935 ;
        RECT 56.325 -147.505 56.810 -138.620 ;
        RECT 63.265 -148.230 63.670 -136.185 ;
        RECT 65.340 -146.330 65.730 -134.905 ;
        RECT 68.500 -142.490 68.855 -131.405 ;
        RECT 72.245 -132.765 72.535 -130.705 ;
        RECT 75.015 -132.165 75.515 -129.115 ;
        RECT 79.985 -132.255 80.395 -129.160 ;
        RECT 79.025 -133.915 79.335 -133.885 ;
        RECT 69.825 -137.635 70.295 -134.645 ;
        RECT 72.175 -140.620 72.490 -138.250 ;
        RECT 73.795 -138.575 74.215 -134.610 ;
        RECT 70.460 -143.330 70.840 -141.955 ;
        RECT 72.900 -144.360 73.245 -141.900 ;
        RECT 74.535 -142.680 74.860 -139.915 ;
        RECT 75.520 -140.645 75.925 -137.315 ;
        RECT 79.025 -140.015 79.340 -133.915 ;
        RECT 80.170 -143.620 80.540 -134.520 ;
        RECT 81.115 -142.555 81.405 -130.720 ;
        RECT 84.565 -132.280 84.975 -129.185 ;
        RECT 89.020 -132.825 89.330 -130.310 ;
        RECT 93.270 -131.125 93.650 -130.745 ;
        RECT 95.400 -131.125 95.780 -130.745 ;
        RECT 82.010 -140.060 82.340 -133.865 ;
        RECT 84.915 -140.590 85.370 -137.315 ;
        RECT 87.275 -138.575 87.820 -134.635 ;
        RECT 91.330 -137.635 91.765 -134.625 ;
        RECT 86.470 -142.680 86.795 -139.915 ;
        RECT 88.985 -140.585 89.400 -138.195 ;
        RECT 92.525 -142.010 92.855 -131.315 ;
        RECT 93.960 -137.675 94.345 -131.890 ;
        RECT 90.715 -143.415 91.050 -142.065 ;
        RECT 94.320 -142.430 94.745 -138.155 ;
        RECT 96.020 -140.665 96.320 -133.625 ;
        RECT 97.140 -141.270 97.440 -134.340 ;
        RECT 98.450 -140.670 98.750 -134.320 ;
        RECT 92.980 -143.340 93.360 -142.960 ;
        RECT 95.175 -143.355 95.555 -142.975 ;
        RECT 99.045 -143.415 99.335 -133.635 ;
        RECT 99.765 -140.640 100.060 -133.815 ;
        RECT 100.895 -141.180 101.195 -134.370 ;
        RECT 101.685 -140.585 101.995 -130.545 ;
        RECT 110.875 -132.300 111.255 -131.920 ;
        RECT 102.480 -140.655 102.780 -133.825 ;
        RECT 103.605 -141.270 103.905 -134.330 ;
        RECT 105.055 -141.395 105.335 -138.360 ;
        RECT 105.815 -140.695 106.095 -134.335 ;
        RECT 106.665 -140.695 106.965 -133.875 ;
        RECT 107.805 -141.440 108.105 -134.285 ;
        RECT 108.450 -137.250 108.830 -136.870 ;
        RECT 108.450 -139.305 108.830 -138.925 ;
        RECT 110.300 -139.425 110.615 -135.100 ;
        RECT 110.910 -137.350 111.190 -135.820 ;
        RECT 111.480 -140.665 111.780 -133.625 ;
        RECT 113.255 -139.910 113.555 -135.850 ;
        RECT 110.775 -142.475 111.155 -142.095 ;
        RECT 114.505 -142.880 114.795 -133.635 ;
        RECT 116.355 -141.180 116.655 -134.370 ;
        RECT 117.145 -140.585 117.455 -131.850 ;
        RECT 117.940 -140.655 118.240 -133.825 ;
        RECT 119.745 -139.925 120.025 -135.835 ;
        RECT 120.515 -141.395 120.795 -138.360 ;
        RECT 123.265 -141.440 123.565 -134.285 ;
        RECT 125.605 -135.670 125.980 -127.470 ;
        RECT 127.350 -136.475 127.650 -125.480 ;
        RECT -1.115 -160.925 -0.815 -153.995 ;
        RECT 0.195 -160.325 0.495 -153.975 ;
        RECT 1.510 -160.295 1.805 -153.470 ;
        RECT 5.350 -160.925 5.650 -153.985 ;
        RECT 7.560 -160.350 7.865 -153.990 ;
        RECT 8.410 -160.350 8.710 -153.530 ;
        RECT 10.220 -156.905 10.600 -156.525 ;
        RECT 12.005 -158.325 12.325 -156.195 ;
        RECT 10.435 -161.615 10.815 -158.595 ;
        RECT 12.615 -159.165 12.895 -156.760 ;
        RECT 13.225 -160.320 13.525 -153.280 ;
        RECT 14.345 -160.925 14.645 -153.995 ;
        RECT 15.655 -160.325 15.955 -153.975 ;
        RECT 16.250 -158.450 16.575 -153.290 ;
        RECT 16.970 -160.295 17.265 -153.470 ;
        RECT 18.100 -160.835 18.400 -154.025 ;
        RECT 18.890 -160.240 19.200 -154.050 ;
        RECT 19.685 -160.310 19.985 -153.480 ;
        RECT 20.810 -160.925 21.110 -153.985 ;
        RECT 22.260 -161.050 22.540 -158.015 ;
        RECT 23.020 -160.350 23.340 -153.990 ;
        RECT 23.870 -160.350 24.170 -153.530 ;
        RECT 25.010 -161.095 25.310 -153.940 ;
        RECT 25.645 -158.950 26.025 -158.570 ;
        RECT 26.350 -163.065 26.710 -156.505 ;
        RECT 27.490 -158.315 27.815 -156.450 ;
        RECT 28.155 -161.660 28.615 -156.975 ;
        RECT 28.940 -159.115 29.390 -150.295 ;
        RECT 31.125 -157.290 31.555 -154.300 ;
        RECT 28.870 -163.005 29.250 -162.625 ;
        RECT 31.760 -162.985 32.140 -161.610 ;
        RECT 32.530 -162.165 32.845 -151.115 ;
        RECT 33.545 -152.420 33.835 -150.360 ;
        RECT 36.330 -151.820 36.805 -148.770 ;
        RECT 41.285 -151.910 41.695 -148.815 ;
        RECT 33.465 -160.275 33.790 -157.905 ;
        RECT 35.115 -158.230 35.515 -154.265 ;
        RECT 34.200 -164.015 34.545 -161.555 ;
        RECT 35.835 -162.335 36.160 -159.570 ;
        RECT 36.820 -160.300 37.225 -156.970 ;
        RECT 41.470 -163.275 41.840 -154.175 ;
        RECT 42.415 -162.210 42.705 -150.375 ;
        RECT 45.865 -151.935 46.275 -148.840 ;
        RECT 50.320 -152.480 50.630 -149.965 ;
        RECT 46.230 -160.245 46.670 -156.970 ;
        RECT 48.610 -158.230 49.135 -154.290 ;
        RECT 47.770 -162.335 48.095 -159.570 ;
        RECT 50.285 -160.240 50.700 -157.850 ;
        RECT 51.315 -161.680 51.630 -150.995 ;
        RECT 52.645 -157.290 53.130 -154.280 ;
        RECT 59.105 -155.370 62.430 -154.780 ;
        RECT 59.105 -155.985 59.855 -155.370 ;
        RECT 61.010 -158.825 61.680 -156.175 ;
        RECT 52.015 -163.070 52.350 -161.720 ;
        RECT 62.970 -174.980 63.420 -155.940 ;
        RECT 64.760 -175.755 65.175 -154.575 ;
        RECT 68.500 -162.155 68.855 -151.070 ;
        RECT 72.245 -152.430 72.535 -150.370 ;
        RECT 75.015 -151.830 75.515 -148.780 ;
        RECT 79.985 -151.920 80.395 -148.825 ;
        RECT 79.025 -153.580 79.335 -153.550 ;
        RECT 69.825 -157.300 70.295 -154.310 ;
        RECT 72.175 -160.285 72.490 -157.915 ;
        RECT 73.795 -158.240 74.215 -154.275 ;
        RECT 70.460 -162.995 70.840 -161.620 ;
        RECT 72.900 -164.025 73.245 -161.565 ;
        RECT 74.535 -162.345 74.860 -159.580 ;
        RECT 75.520 -160.310 75.925 -156.980 ;
        RECT 79.025 -159.680 79.340 -153.580 ;
        RECT 80.170 -163.285 80.540 -154.185 ;
        RECT 81.115 -162.220 81.405 -150.385 ;
        RECT 84.565 -151.945 84.975 -148.850 ;
        RECT 89.020 -152.490 89.330 -149.975 ;
        RECT 93.270 -150.790 93.650 -150.410 ;
        RECT 95.400 -150.790 95.780 -150.410 ;
        RECT 82.010 -159.725 82.340 -153.530 ;
        RECT 84.915 -160.255 85.370 -156.980 ;
        RECT 87.275 -158.240 87.820 -154.300 ;
        RECT 91.330 -157.300 91.765 -154.290 ;
        RECT 86.470 -162.345 86.795 -159.580 ;
        RECT 88.985 -160.250 89.400 -157.860 ;
        RECT 92.525 -161.675 92.855 -150.980 ;
        RECT 93.960 -157.340 94.345 -151.555 ;
        RECT 90.715 -163.080 91.050 -161.730 ;
        RECT 94.320 -162.095 94.745 -157.820 ;
        RECT 96.020 -160.330 96.320 -153.290 ;
        RECT 97.140 -160.935 97.440 -154.005 ;
        RECT 98.450 -160.335 98.750 -153.985 ;
        RECT 92.980 -163.005 93.360 -162.625 ;
        RECT 95.175 -163.020 95.555 -162.640 ;
        RECT 99.045 -163.080 99.335 -153.300 ;
        RECT 99.765 -160.305 100.060 -153.480 ;
        RECT 100.895 -160.845 101.195 -154.035 ;
        RECT 101.685 -160.250 101.995 -150.210 ;
        RECT 110.875 -151.965 111.255 -151.585 ;
        RECT 102.480 -160.320 102.780 -153.490 ;
        RECT 103.605 -160.935 103.905 -153.995 ;
        RECT 105.055 -161.060 105.335 -158.025 ;
        RECT 105.815 -160.360 106.095 -154.000 ;
        RECT 106.665 -160.360 106.965 -153.540 ;
        RECT 107.805 -161.105 108.105 -153.950 ;
        RECT 108.450 -156.915 108.830 -156.535 ;
        RECT 108.450 -158.970 108.830 -158.590 ;
        RECT 110.300 -159.090 110.615 -154.765 ;
        RECT 110.910 -157.015 111.190 -155.485 ;
        RECT 111.480 -160.330 111.780 -153.290 ;
        RECT 113.255 -159.575 113.555 -155.515 ;
        RECT 110.775 -162.140 111.155 -161.760 ;
        RECT 114.505 -162.545 114.795 -153.300 ;
        RECT 116.355 -160.845 116.655 -154.035 ;
        RECT 117.145 -160.250 117.455 -151.515 ;
        RECT 117.940 -160.320 118.240 -153.490 ;
        RECT 119.745 -159.590 120.025 -155.500 ;
        RECT 120.515 -161.060 120.795 -158.025 ;
        RECT 123.265 -161.105 123.565 -153.950 ;
        RECT 125.190 -155.185 125.565 -147.345 ;
        RECT 127.045 -155.935 127.345 -145.395 ;
        RECT 67.400 -180.065 67.700 -173.025 ;
        RECT 69.175 -179.310 69.475 -175.250 ;
        RECT 70.425 -178.195 70.745 -173.035 ;
        RECT 72.275 -180.580 72.575 -173.770 ;
        RECT 73.065 -179.985 73.375 -173.795 ;
        RECT 73.860 -180.055 74.160 -173.225 ;
        RECT 75.665 -179.325 75.945 -175.235 ;
        RECT 76.435 -180.795 76.715 -177.760 ;
        RECT 79.185 -180.840 79.485 -173.685 ;
      LAYER Metal3 ;
        RECT 93.225 145.560 95.820 145.990 ;
        RECT 93.905 144.435 111.275 144.775 ;
        RECT 10.280 139.545 28.005 139.865 ;
        RECT 108.430 139.465 111.275 139.845 ;
        RECT -8.205 138.170 12.500 138.465 ;
        RECT -8.385 137.305 13.085 137.600 ;
        RECT 25.695 137.425 29.595 137.910 ;
        RECT 108.405 137.390 110.690 137.815 ;
        RECT 10.445 134.770 28.745 135.155 ;
        RECT 94.160 134.235 111.345 134.720 ;
        RECT 26.325 133.450 29.390 133.775 ;
        RECT 92.970 133.320 95.565 133.770 ;
        RECT -8.245 130.695 55.635 131.115 ;
        RECT 64.310 130.820 127.755 131.440 ;
        RECT -6.605 129.150 56.835 129.640 ;
        RECT 62.215 128.865 125.940 129.435 ;
        RECT 93.025 125.835 95.620 126.265 ;
        RECT 93.705 124.710 111.075 125.050 ;
        RECT 10.235 119.855 27.960 120.175 ;
        RECT 108.230 119.740 111.075 120.120 ;
        RECT -8.250 118.480 12.455 118.775 ;
        RECT -8.430 117.615 13.040 117.910 ;
        RECT 25.650 117.735 29.550 118.220 ;
        RECT 108.205 117.665 110.490 118.090 ;
        RECT 10.400 115.080 28.700 115.465 ;
        RECT 93.960 114.510 111.145 114.995 ;
        RECT 26.280 113.760 29.345 114.085 ;
        RECT 92.770 113.595 95.365 114.045 ;
        RECT -8.245 111.195 55.635 111.615 ;
        RECT 64.610 111.070 128.055 111.690 ;
        RECT -6.605 109.650 56.835 110.140 ;
        RECT 62.515 109.115 126.240 109.685 ;
        RECT 93.180 106.190 95.775 106.620 ;
        RECT 93.860 105.065 111.230 105.405 ;
        RECT 10.425 100.145 28.150 100.465 ;
        RECT 108.385 100.095 111.230 100.475 ;
        RECT -8.060 98.770 12.645 99.065 ;
        RECT -8.240 97.905 13.230 98.200 ;
        RECT 25.840 98.025 29.740 98.510 ;
        RECT 108.360 98.020 110.645 98.445 ;
        RECT 10.590 95.370 28.890 95.755 ;
        RECT 94.115 94.865 111.300 95.350 ;
        RECT 26.470 94.050 29.535 94.375 ;
        RECT 92.925 93.950 95.520 94.400 ;
        RECT -8.035 91.155 55.845 91.575 ;
        RECT 64.630 91.410 128.075 92.030 ;
        RECT -6.395 89.610 57.045 90.100 ;
        RECT 62.535 89.455 126.260 90.025 ;
        RECT 93.180 86.395 95.775 86.825 ;
        RECT 93.860 85.270 111.230 85.610 ;
        RECT 10.230 80.305 27.955 80.625 ;
        RECT 108.385 80.300 111.230 80.680 ;
        RECT -8.255 78.930 12.450 79.225 ;
        RECT -8.435 78.065 13.035 78.360 ;
        RECT 25.645 78.185 29.545 78.670 ;
        RECT 108.360 78.225 110.645 78.650 ;
        RECT 10.395 75.530 28.695 75.915 ;
        RECT 94.115 75.070 111.300 75.555 ;
        RECT 26.275 74.210 29.340 74.535 ;
        RECT 92.925 74.155 95.520 74.605 ;
        RECT -8.080 71.365 55.800 71.785 ;
        RECT 64.630 71.675 128.075 72.295 ;
        RECT -6.440 69.820 57.000 70.310 ;
        RECT 62.535 69.720 126.260 70.290 ;
        RECT 93.100 66.640 95.695 67.070 ;
        RECT 93.780 65.515 111.150 65.855 ;
        RECT 10.100 60.595 27.825 60.915 ;
        RECT 108.305 60.545 111.150 60.925 ;
        RECT -8.385 59.220 12.320 59.515 ;
        RECT -8.565 58.355 12.905 58.650 ;
        RECT 25.515 58.475 29.415 58.960 ;
        RECT 108.280 58.470 110.565 58.895 ;
        RECT 10.265 55.820 28.565 56.205 ;
        RECT 94.035 55.315 111.220 55.800 ;
        RECT 26.145 54.500 29.210 54.825 ;
        RECT 92.845 54.400 95.440 54.850 ;
        RECT -8.385 51.735 55.495 52.155 ;
        RECT 64.530 51.970 127.975 52.590 ;
        RECT -6.745 50.190 56.695 50.680 ;
        RECT 62.435 50.015 126.160 50.585 ;
        RECT 93.205 46.925 95.800 47.355 ;
        RECT 93.885 45.800 111.255 46.140 ;
        RECT 10.230 40.835 27.955 41.155 ;
        RECT 108.410 40.830 111.255 41.210 ;
        RECT -8.255 39.460 12.450 39.755 ;
        RECT -8.435 38.595 13.035 38.890 ;
        RECT 25.645 38.715 29.545 39.200 ;
        RECT 108.385 38.755 110.670 39.180 ;
        RECT 10.395 36.060 28.695 36.445 ;
        RECT 94.140 35.600 111.325 36.085 ;
        RECT 26.275 34.740 29.340 35.065 ;
        RECT 92.950 34.685 95.545 35.135 ;
        RECT -8.290 31.960 55.590 32.380 ;
        RECT 64.790 31.815 128.235 32.435 ;
        RECT -6.650 30.415 56.790 30.905 ;
        RECT 62.695 29.860 126.420 30.430 ;
        RECT 93.205 26.955 95.800 27.385 ;
        RECT 93.885 25.830 111.255 26.170 ;
        RECT 10.180 21.025 27.905 21.345 ;
        RECT 108.410 20.860 111.255 21.240 ;
        RECT -8.305 19.650 12.400 19.945 ;
        RECT -8.485 18.785 12.985 19.080 ;
        RECT 25.595 18.905 29.495 19.390 ;
        RECT 108.385 18.785 110.670 19.210 ;
        RECT 10.345 16.250 28.645 16.635 ;
        RECT 94.140 15.630 111.325 16.115 ;
        RECT 26.225 14.930 29.290 15.255 ;
        RECT 92.950 14.715 95.545 15.165 ;
        RECT -8.290 12.150 55.590 12.570 ;
        RECT 64.900 11.925 128.345 12.545 ;
        RECT -6.650 10.605 56.790 11.095 ;
        RECT 62.805 9.970 126.530 10.540 ;
        RECT 93.205 7.290 95.800 7.720 ;
        RECT 93.885 6.165 111.255 6.505 ;
        RECT 10.150 1.230 27.875 1.550 ;
        RECT 108.410 1.195 111.255 1.575 ;
        RECT -8.335 -0.145 12.370 0.150 ;
        RECT -8.515 -1.010 12.955 -0.715 ;
        RECT 25.565 -0.890 29.465 -0.405 ;
        RECT 108.385 -0.880 110.670 -0.455 ;
        RECT 10.315 -3.545 28.615 -3.160 ;
        RECT 94.140 -4.035 111.325 -3.550 ;
        RECT 26.195 -4.865 29.260 -4.540 ;
        RECT 92.950 -4.950 95.545 -4.500 ;
        RECT -8.450 -8.035 56.200 -7.550 ;
        RECT 64.270 -7.765 128.055 -7.135 ;
        RECT -6.505 -9.410 57.905 -8.870 ;
        RECT 62.340 -9.060 126.325 -8.525 ;
        RECT 93.245 -12.550 95.840 -12.120 ;
        RECT 93.925 -13.675 111.295 -13.335 ;
        RECT 10.300 -18.565 28.025 -18.245 ;
        RECT 108.450 -18.645 111.295 -18.265 ;
        RECT -8.185 -19.940 12.520 -19.645 ;
        RECT -8.365 -20.805 13.105 -20.510 ;
        RECT 25.715 -20.685 29.615 -20.200 ;
        RECT 108.425 -20.720 110.710 -20.295 ;
        RECT 10.465 -23.340 28.765 -22.955 ;
        RECT 94.180 -23.875 111.365 -23.390 ;
        RECT 26.345 -24.660 29.410 -24.335 ;
        RECT 92.990 -24.790 95.585 -24.340 ;
        RECT -8.225 -27.415 55.655 -26.995 ;
        RECT 64.330 -27.290 127.775 -26.670 ;
        RECT -6.585 -28.960 56.855 -28.470 ;
        RECT 62.235 -29.245 125.960 -28.675 ;
        RECT 93.045 -32.275 95.640 -31.845 ;
        RECT 93.725 -33.400 111.095 -33.060 ;
        RECT 10.255 -38.255 27.980 -37.935 ;
        RECT 108.250 -38.370 111.095 -37.990 ;
        RECT -8.230 -39.630 12.475 -39.335 ;
        RECT -8.410 -40.495 13.060 -40.200 ;
        RECT 25.670 -40.375 29.570 -39.890 ;
        RECT 108.225 -40.445 110.510 -40.020 ;
        RECT 10.420 -43.030 28.720 -42.645 ;
        RECT 93.980 -43.600 111.165 -43.115 ;
        RECT 26.300 -44.350 29.365 -44.025 ;
        RECT 92.790 -44.515 95.385 -44.065 ;
        RECT -8.225 -46.915 55.655 -46.495 ;
        RECT 64.630 -47.040 128.075 -46.420 ;
        RECT -6.585 -48.460 56.855 -47.970 ;
        RECT 62.535 -48.995 126.260 -48.425 ;
        RECT 93.200 -51.920 95.795 -51.490 ;
        RECT 93.880 -53.045 111.250 -52.705 ;
        RECT 10.445 -57.965 28.170 -57.645 ;
        RECT 108.405 -58.015 111.250 -57.635 ;
        RECT -8.040 -59.340 12.665 -59.045 ;
        RECT -8.220 -60.205 13.250 -59.910 ;
        RECT 25.860 -60.085 29.760 -59.600 ;
        RECT 108.380 -60.090 110.665 -59.665 ;
        RECT 10.610 -62.740 28.910 -62.355 ;
        RECT 94.135 -63.245 111.320 -62.760 ;
        RECT 26.490 -64.060 29.555 -63.735 ;
        RECT 92.945 -64.160 95.540 -63.710 ;
        RECT -8.015 -66.955 55.865 -66.535 ;
        RECT 64.650 -66.700 128.095 -66.080 ;
        RECT -6.375 -68.500 57.065 -68.010 ;
        RECT 62.555 -68.655 126.280 -68.085 ;
        RECT 93.200 -71.715 95.795 -71.285 ;
        RECT 93.880 -72.840 111.250 -72.500 ;
        RECT 10.250 -77.805 27.975 -77.485 ;
        RECT 108.405 -77.810 111.250 -77.430 ;
        RECT -8.235 -79.180 12.470 -78.885 ;
        RECT -8.415 -80.045 13.055 -79.750 ;
        RECT 25.665 -79.925 29.565 -79.440 ;
        RECT 108.380 -79.885 110.665 -79.460 ;
        RECT 10.415 -82.580 28.715 -82.195 ;
        RECT 94.135 -83.040 111.320 -82.555 ;
        RECT 26.295 -83.900 29.360 -83.575 ;
        RECT 92.945 -83.955 95.540 -83.505 ;
        RECT -8.060 -86.745 55.820 -86.325 ;
        RECT 64.650 -86.435 128.095 -85.815 ;
        RECT -6.420 -88.290 57.020 -87.800 ;
        RECT 62.555 -88.390 126.280 -87.820 ;
        RECT 93.120 -91.470 95.715 -91.040 ;
        RECT 93.800 -92.595 111.170 -92.255 ;
        RECT 10.120 -97.515 27.845 -97.195 ;
        RECT 108.325 -97.565 111.170 -97.185 ;
        RECT -8.365 -98.890 12.340 -98.595 ;
        RECT -8.545 -99.755 12.925 -99.460 ;
        RECT 25.535 -99.635 29.435 -99.150 ;
        RECT 108.300 -99.640 110.585 -99.215 ;
        RECT 10.285 -102.290 28.585 -101.905 ;
        RECT 94.055 -102.795 111.240 -102.310 ;
        RECT 26.165 -103.610 29.230 -103.285 ;
        RECT 92.865 -103.710 95.460 -103.260 ;
        RECT -8.365 -106.375 55.515 -105.955 ;
        RECT 64.550 -106.140 127.995 -105.520 ;
        RECT -6.725 -107.920 56.715 -107.430 ;
        RECT 62.455 -108.095 126.180 -107.525 ;
        RECT 93.225 -111.185 95.820 -110.755 ;
        RECT 93.905 -112.310 111.275 -111.970 ;
        RECT 10.250 -117.275 27.975 -116.955 ;
        RECT 108.430 -117.280 111.275 -116.900 ;
        RECT -8.235 -118.650 12.470 -118.355 ;
        RECT -8.415 -119.515 13.055 -119.220 ;
        RECT 25.665 -119.395 29.565 -118.910 ;
        RECT 108.405 -119.355 110.690 -118.930 ;
        RECT 10.415 -122.050 28.715 -121.665 ;
        RECT 94.160 -122.510 111.345 -122.025 ;
        RECT 26.295 -123.370 29.360 -123.045 ;
        RECT 92.970 -123.425 95.565 -122.975 ;
        RECT -8.270 -126.150 55.610 -125.730 ;
        RECT 64.810 -126.295 128.255 -125.675 ;
        RECT -6.630 -127.695 56.810 -127.205 ;
        RECT 62.715 -128.250 126.440 -127.680 ;
        RECT 93.225 -131.155 95.820 -130.725 ;
        RECT 93.905 -132.280 111.275 -131.940 ;
        RECT 10.200 -137.085 27.925 -136.765 ;
        RECT 108.430 -137.250 111.275 -136.870 ;
        RECT -8.285 -138.460 12.420 -138.165 ;
        RECT -8.465 -139.325 13.005 -139.030 ;
        RECT 25.615 -139.205 29.515 -138.720 ;
        RECT 108.405 -139.325 110.690 -138.900 ;
        RECT 10.365 -141.860 28.665 -141.475 ;
        RECT 94.160 -142.480 111.345 -141.995 ;
        RECT 26.245 -143.180 29.310 -142.855 ;
        RECT 92.970 -143.395 95.565 -142.945 ;
        RECT -8.270 -145.960 55.610 -145.540 ;
        RECT 64.920 -146.185 128.365 -145.565 ;
        RECT -6.630 -147.505 56.810 -147.015 ;
        RECT 62.825 -148.140 126.550 -147.570 ;
        RECT 93.225 -150.820 95.820 -150.390 ;
        RECT 93.905 -151.945 111.275 -151.605 ;
        RECT 10.170 -156.880 27.895 -156.560 ;
        RECT 108.430 -156.915 111.275 -156.535 ;
        RECT -8.315 -158.255 12.390 -157.960 ;
        RECT -8.495 -159.120 12.975 -158.825 ;
        RECT 25.585 -159.000 29.485 -158.515 ;
        RECT 108.405 -158.990 110.690 -158.565 ;
        RECT 10.335 -161.655 28.635 -161.270 ;
        RECT 94.160 -162.145 111.345 -161.660 ;
        RECT 26.215 -162.975 29.280 -162.650 ;
        RECT 92.970 -163.060 95.565 -162.610 ;
  END
END fa16b_rev
END LIBRARY

